* SPICE NETLIST
***************************************

.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT WELLTAP
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6
** N=7 EP=6 IP=0 FDC=4
M0 7 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 7 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 11 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 10 A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 10 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7
** N=9 EP=7 IP=0 FDC=6
M0 ZN B2 8 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 8 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 8 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_6
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS
** N=10 EP=7 IP=0 FDC=8
M0 9 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 8 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 8 A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MUX2_X1 A S B VSS VDD Z 7
** N=13 EP=7 IP=0 FDC=12
M0 VSS S 8 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 12 A VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 9 8 12 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 13 S 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=715 $Y=90 $D=1
M4 VSS B 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=905 $Y=90 $D=1
M5 Z 9 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 VDD S 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M7 10 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M8 9 S 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M9 11 8 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=715 $Y=995 $D=0
M10 VDD B 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=905 $Y=995 $D=0
M11 Z 9 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6
** N=10 EP=6 IP=0 FDC=10
M0 10 A 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 10 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 8 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 8 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 7 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 9 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_11
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=12
X1 3 4 5 1 2 6 1 MUX2_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7
** N=13 EP=7 IP=0 FDC=16
M0 12 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 12 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 9 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 9 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 13 A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 10 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 8 A S VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 9 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 9 A 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 10 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 10 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN C2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 8 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 10 A 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6
** N=7 EP=6 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 7 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN 6
** N=8 EP=6 IP=0 FDC=6
M0 7 A1 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8
** N=20 EP=8 IP=0 FDC=28
M0 VSS 9 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 18 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 9 A 18 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 10 CI 9 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 10 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 12 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 12 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 14 9 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 19 CI 14 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 20 B 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 14 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 9 CO VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 15 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 9 A 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 11 CI 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 13 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 13 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 14 9 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 16 CI 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 17 B 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 17 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 14 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 7 A1 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 6 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 8 A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_24
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=3 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT AOI222_X1 C2 C1 VDD B1 B2 A2 VSS A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=1.2035e-13 AS=5.81e-14 PD=1.41e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 13 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=1.2035e-13 PD=1.11e-06 PS=1.41e-06 $X=675 $Y=90 $D=1
M3 VSS B2 13 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=865 $Y=90 $D=1
M4 14 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1055 $Y=90 $D=1
M5 ZN A1 14 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1245 $Y=90 $D=1
M6 10 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M7 VDD C1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M8 10 B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=675 $Y=680 $D=0
M9 11 B2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=865 $Y=680 $D=0
M10 ZN A2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1055 $Y=680 $D=0
M11 11 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1245 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=6
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD
** N=10 EP=7 IP=0 FDC=8
M0 VSS B2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 8 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 8 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 10 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT OAI222_X1 C2 C1 VSS B1 B2 A2 VDD A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 10 B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=710 $Y=90 $D=1
M3 11 B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=900 $Y=90 $D=1
M4 ZN A2 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1090 $Y=90 $D=1
M5 11 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1280 $Y=90 $D=1
M6 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M7 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M8 13 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=710 $Y=680 $D=0
M9 VDD B2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=900 $Y=680 $D=0
M10 14 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1090 $Y=680 $D=0
M11 ZN A1 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1280 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 9 A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X2 A1 ZN A2 A3 VSS VDD
** N=10 EP=6 IP=0 FDC=12
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M7 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M8 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M9 9 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M10 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M11 VDD A3 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6
** N=10 EP=6 IP=0 FDC=10
M0 7 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 10 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 10 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 9 A 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 8 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 8 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 5 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X2 A VDD B1 ZN B2 VSS
** N=9 EP=6 IP=0 FDC=12
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M7 7 A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M8 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M9 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M10 ZN B1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M11 7 B2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=10
X1 2 3 4 5 1 1 XOR2_X1 $T=1140 0 0 0 $X=1025 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_34
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN 7
** N=10 EP=7 IP=0 FDC=8
M0 VSS A1 8 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 8 A2 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 8 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 8 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 9 A1 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 10 A2 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=24
X0 1 2 3 4 5 6 11 MUX2_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 7 8 9 4 5 10 11 MUX2_X1 $T=1330 0 0 0 $X=1215 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=11 FDC=16
X0 1 2 3 4 5 AND2_X1 $T=1140 0 0 0 $X=1025 $Y=-115
X1 4 6 7 8 3 3 XOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5 6 7
** N=7 EP=7 IP=13 FDC=18
X0 1 2 3 4 5 6 7 AOI22_X1 $T=1140 0 0 0 $X=1025 $Y=-115
X1 3 2 4 1 7 7 XOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=13 FDC=22
X0 1 2 3 4 5 6 4 MUX2_X1 $T=1140 0 0 0 $X=1025 $Y=-115
X1 5 7 8 9 4 4 XOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6
** N=6 EP=6 IP=9 FDC=12
X1 3 4 5 1 2 6 1 MUX2_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT floatingadder a[2] a[10] a[16] b[5] b[4] b[3] a[6] b[2] b[10] b[16] a[5] a[4] a[3] b[6] b[15] b[14] a[12] a[11] a[1] a[9]
+ a[8] a[7] a[15] a[14] b[12] b[11] b[1] b[9] b[8] b[7] a[17] b[17] b[13] a[0] a[13] b[0] b[28] b[30] a[30] b[27]
+ b[23] b[24] b[26] a[24] a[23] b[25] a[25] a[28] a[19] b[18] b[19] a[18] a[22] b[29] a[29] b[21] a[21] b[22] a[20] b[20]
+ a[31] b[31] sum[30] a[27] a[26] VSS VDD sum[31] sum[29] sum[20] sum[26] sum[2] sum[22] sum[23] sum[5] sum[21] sum[11] sum[25] sum[14] sum[10]
+ sum[3] sum[16] sum[18] sum[17] sum[15] sum[13] sum[9] sum[8] sum[12] sum[24] sum[28] sum[1] sum[0] sum[6] sum[27] sum[7] sum[19] sum[4] carry clk
** N=975 EP=100 IP=13304 FDC=7024
M0 VSS 492 493 VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=3045 $Y=11915 $D=1
M1 18 493 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=3235 $Y=11915 $D=1
M2 VSS 493 18 VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=3425 $Y=11915 $D=1
M3 494 495 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=4575 $Y=9490 $D=1
M4 VSS 495 494 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=4765 $Y=9490 $D=1
M5 968 499 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=4955 $Y=9490 $D=1
M6 495 497 968 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=5145 $Y=9490 $D=1
M7 494 497 68 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=5530 $Y=9490 $D=1
M8 68 497 494 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=5720 $Y=9490 $D=1
M9 494 499 68 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=5910 $Y=9490 $D=1
M10 68 499 494 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=6100 $Y=9490 $D=1
M11 503 109 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=11055 $Y=8895 $D=1
M12 VSS 502 503 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=11245 $Y=8895 $D=1
M13 74 503 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=11435 $Y=8895 $D=1
M14 969 109 74 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=11625 $Y=8895 $D=1
M15 VSS 502 969 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=11815 $Y=8895 $D=1
M16 970 502 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=12005 $Y=8895 $D=1
M17 74 109 970 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=12195 $Y=8895 $D=1
M18 VSS 503 74 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=12385 $Y=8895 $D=1
M19 971 366 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=33270 $Y=12290 $D=1
M20 318 516 971 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33460 $Y=12290 $D=1
M21 972 516 318 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33650 $Y=12290 $D=1
M22 VSS 366 972 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=33840 $Y=12290 $D=1
M23 523 519 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=35350 $Y=31890 $D=1
M24 VSS 518 523 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=35540 $Y=31890 $D=1
M25 523 518 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=35730 $Y=31890 $D=1
M26 VSS 519 523 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=7.2625e-14 AS=5.81e-14 PD=1.18e-06 PS=1.11e-06 $X=35920 $Y=31890 $D=1
M27 973 524 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=7.2625e-14 PD=1.11e-06 PS=1.18e-06 $X=36145 $Y=31890 $D=1
M28 526 343 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=36295 $Y=42700 $D=1
M29 523 520 973 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=36335 $Y=31890 $D=1
M30 VSS 375 526 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=36485 $Y=42700 $D=1
M31 974 520 523 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=36525 $Y=31890 $D=1
M32 526 378 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=36675 $Y=42700 $D=1
M33 VSS 524 974 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=36715 $Y=31890 $D=1
M34 VSS 382 526 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=36865 $Y=42700 $D=1
M35 363 526 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=37055 $Y=42495 $D=1
M36 VDD 492 493 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=3045 $Y=10890 $D=0
M37 18 493 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3235 $Y=10890 $D=0
M38 VDD 493 18 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3425 $Y=10890 $D=0
M39 68 495 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=4575 $Y=10080 $D=0
M40 VDD 495 68 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4765 $Y=10080 $D=0
M41 495 499 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4955 $Y=10080 $D=0
M42 VDD 497 495 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=5145 $Y=10080 $D=0
M43 68 497 496 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=5530 $Y=10080 $D=0
M44 961 497 68 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5720 $Y=10080 $D=0
M45 VDD 499 961 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5910 $Y=10080 $D=0
M46 496 499 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=6100 $Y=10080 $D=0
M47 962 109 503 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=11055 $Y=8090 $D=0
M48 VDD 502 962 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=11245 $Y=8090 $D=0
M49 501 503 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=11435 $Y=8090 $D=0
M50 74 109 501 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=11625 $Y=8090 $D=0
M51 501 502 74 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=11815 $Y=8090 $D=0
M52 74 502 501 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=12005 $Y=8090 $D=0
M53 501 109 74 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=12195 $Y=8090 $D=0
M54 VDD 503 501 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=12385 $Y=8090 $D=0
M55 318 366 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=33270 $Y=12880 $D=0
M56 VDD 516 318 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33460 $Y=12880 $D=0
M57 318 516 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33650 $Y=12880 $D=0
M58 VDD 366 318 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=33840 $Y=12880 $D=0
M59 963 519 525 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=35350 $Y=32480 $D=0
M60 VDD 518 963 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35540 $Y=32480 $D=0
M61 964 518 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35730 $Y=32480 $D=0
M62 525 519 964 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=1.1025e-13 AS=8.82e-14 PD=1.61e-06 PS=1.54e-06 $X=35920 $Y=32480 $D=0
M63 523 524 525 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.1025e-13 PD=1.54e-06 PS=1.61e-06 $X=36145 $Y=32480 $D=0
M64 965 343 526 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=36295 $Y=41690 $D=0
M65 525 520 523 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=36335 $Y=32480 $D=0
M66 966 375 965 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=36485 $Y=41690 $D=0
M67 523 520 525 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=36525 $Y=32480 $D=0
M68 967 378 966 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=36675 $Y=41690 $D=0
M69 525 524 523 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=36715 $Y=32480 $D=0
M70 VDD 382 967 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=36865 $Y=41690 $D=0
M71 363 526 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=37055 $Y=41690 $D=0
X5706 43 VSS 498 121 VDD VSS NAND2_X1 $T=4990 15000 0 0 $X=4875 $Y=14885
X5707 61 VSS 68 544 VDD VSS NAND2_X1 $T=5940 17800 1 0 $X=5825 $Y=16285
X5708 547 VSS 60 65 VDD VSS NAND2_X1 $T=7080 17800 0 0 $X=6965 $Y=17685
X5709 731 VSS 854 72 VDD VSS NAND2_X1 $T=7650 23400 0 180 $X=6965 $Y=21885
X5710 949 VSS 83 577 VDD VSS NAND2_X1 $T=7270 31800 1 0 $X=7155 $Y=30285
X5711 555 VSS 93 730 VDD VSS NAND2_X1 $T=8410 23400 1 180 $X=7725 $Y=23285
X5712 856 VSS 499 553 VDD VSS NAND2_X1 $T=8410 9400 0 0 $X=8295 $Y=9285
X5713 556 VSS 59 101 VDD VSS NAND2_X1 $T=9360 12200 1 180 $X=8675 $Y=12085
X5714 557 VSS 554 98 VDD VSS NAND2_X1 $T=9360 17800 1 180 $X=8675 $Y=17685
X5715 547 VSS 140 731 VDD VSS NAND2_X1 $T=8790 20600 0 0 $X=8675 $Y=20485
X5716 547 VSS 110 555 VDD VSS NAND2_X1 $T=8790 23400 1 0 $X=8675 $Y=21885
X5717 547 VSS 118 557 VDD VSS NAND2_X1 $T=9550 17800 1 0 $X=9435 $Y=16285
X5718 741 VSS 574 172 VDD VSS NAND2_X1 $T=11450 12200 0 180 $X=10765 $Y=10685
X5719 569 VSS 741 558 VDD VSS NAND2_X1 $T=12590 12200 1 0 $X=12475 $Y=10685
X5720 741 VSS 111 755 VDD VSS NAND2_X1 $T=13160 12200 1 0 $X=13045 $Y=10685
X5721 559 VSS 569 894 VDD VSS NAND2_X1 $T=14300 12200 0 180 $X=13615 $Y=10685
X5722 111 VSS 559 578 VDD VSS NAND2_X1 $T=13920 12200 0 0 $X=13805 $Y=12085
X5723 156 VSS 108 505 VDD VSS NAND2_X1 $T=14300 23400 1 0 $X=14185 $Y=21885
X5724 579 VSS 186 584 VDD VSS NAND2_X1 $T=16770 17800 0 0 $X=16655 $Y=17685
X5725 862 VSS 213 760 VDD VSS NAND2_X1 $T=19050 29000 0 0 $X=18935 $Y=28885
X5726 763 VSS 863 506 VDD VSS NAND2_X1 $T=19810 20600 1 0 $X=19695 $Y=19085
X5727 597 VSS 223 601 VDD VSS NAND2_X1 $T=21900 6600 1 0 $X=21785 $Y=5085
X5728 783 VSS 270 870 VDD VSS NAND2_X1 $T=25510 37400 1 0 $X=25395 $Y=35885
X5729 790 VSS 304 628 VDD VSS NAND2_X1 $T=27600 26200 1 0 $X=27485 $Y=24685
X5730 644 VSS 641 638 VDD VSS NAND2_X1 $T=30640 3800 0 0 $X=30525 $Y=3685
X5731 139 VSS 638 388 VDD VSS NAND2_X1 $T=31020 12200 0 0 $X=30905 $Y=12085
X5732 644 VSS 647 799 VDD 975 NAND2_X1 $T=32160 1000 0 0 $X=32045 $Y=885
X5733 313 VSS 339 650 VDD VSS NAND2_X1 $T=32350 17800 1 0 $X=32235 $Y=16285
X5734 905 VSS 658 415 VDD VSS NAND2_X1 $T=33870 23400 0 0 $X=33755 $Y=23285
X5735 807 VSS 879 414 VDD VSS NAND2_X1 $T=34060 23400 1 0 $X=33945 $Y=21885
X5736 372 VSS 385 906 VDD VSS NAND2_X1 $T=34630 37400 0 180 $X=33945 $Y=35885
X5737 347 VSS 659 519 VDD VSS NAND2_X1 $T=34250 31800 1 0 $X=34135 $Y=30285
X5738 659 VSS 660 358 VDD VSS NAND2_X1 $T=34440 29000 0 0 $X=34325 $Y=28885
X5739 361 VSS 669 518 VDD VSS NAND2_X1 $T=34630 23400 1 0 $X=34515 $Y=21885
X5740 673 VSS 388 672 VDD VSS NAND2_X1 $T=37480 3800 0 0 $X=37365 $Y=3685
X5741 333 VSS 675 911 VDD VSS NAND2_X1 $T=37670 12200 0 0 $X=37555 $Y=12085
X5742 391 VSS 385 528 VDD VSS NAND2_X1 $T=38810 31800 1 180 $X=38125 $Y=31685
X5743 371 VSS 530 417 VDD VSS NAND2_X1 $T=39570 23400 0 0 $X=39455 $Y=23285
X5744 371 VSS 679 684 VDD VSS NAND2_X1 $T=40140 34600 0 180 $X=39455 $Y=33085
X5745 679 VSS 691 683 VDD VSS NAND2_X1 $T=40330 31800 0 180 $X=39645 $Y=30285
X5746 408 VSS 437 686 VDD VSS NAND2_X1 $T=39950 20600 0 0 $X=39835 $Y=20485
X5747 530 VSS 419 373 VDD VSS NAND2_X1 $T=40140 23400 0 0 $X=40025 $Y=23285
X5748 415 VSS 419 687 VDD VSS NAND2_X1 $T=40140 26200 1 0 $X=40025 $Y=24685
X5749 371 VSS 691 689 VDD VSS NAND2_X1 $T=40330 29000 0 0 $X=40215 $Y=28885
X5750 823 VSS 828 sum[22] VDD VSS NAND2_X1 $T=41280 20600 1 0 $X=41165 $Y=19085
X5751 920 VSS 530 950 VDD VSS NAND2_X1 $T=41280 20600 0 0 $X=41165 $Y=20485
X5752 696 VSS 419 829 VDD VSS NAND2_X1 $T=41850 31800 0 0 $X=41735 $Y=31685
X5753 379 VSS 388 438 VDD VSS NAND2_X1 $T=42230 23400 0 0 $X=42115 $Y=23285
X5754 419 VSS 691 832 VDD VSS NAND2_X1 $T=42800 29000 1 180 $X=42115 $Y=28885
X5755 830 VSS 419 697 VDD VSS NAND2_X1 $T=42230 31800 1 0 $X=42115 $Y=30285
X5756 716 VSS 412 379 VDD VSS NAND2_X1 $T=43370 17800 1 180 $X=42685 $Y=17685
X5757 440 VSS 530 704 VDD VSS NAND2_X1 $T=43750 26200 1 0 $X=43635 $Y=24685
X5758 408 VSS 826 708 VDD VSS NAND2_X1 $T=43750 43000 1 0 $X=43635 $Y=41485
X5759 435 VSS 388 714 VDD VSS NAND2_X1 $T=44700 17800 1 180 $X=44015 $Y=17685
X5760 388 VSS 716 398 VDD VSS NAND2_X1 $T=46030 17800 1 180 $X=45345 $Y=17685
X5761 408 VSS 701 715 VDD VSS NAND2_X1 $T=46220 43000 0 0 $X=46105 $Y=42885
X5762 516 333 366 VSS VDD NOR2_X2 $T=34060 12200 0 0 $X=33945 $Y=12085
X5763 435 429 366 VSS VDD NOR2_X2 $T=45840 17800 1 0 $X=45725 $Y=16285
X5764 366 420 716 VSS VDD NOR2_X2 $T=47170 15000 1 180 $X=46105 $Y=14885
X5790 VDD 111 VDD 55 52 VSS 49 89 AOI221_X1 $T=5940 29000 0 180 $X=4685 $Y=27485
X5791 62 111 VDD 69 72 VSS 68 82 AOI221_X1 $T=5940 29000 1 0 $X=5825 $Y=27485
X5792 52 102 VDD 74 79 VSS 551 549 AOI221_X1 $T=6320 26200 0 0 $X=6205 $Y=26085
X5793 106 52 VDD 95 98 VSS 68 137 AOI221_X1 $T=7650 17800 0 0 $X=7535 $Y=17685
X5794 636 344 VDD 359 351 VSS 336 368 AOI221_X1 $T=34440 26200 0 0 $X=34325 $Y=26085
X5795 351 320 VDD 371 374 VSS 514 814 AOI221_X1 $T=35770 31800 1 0 $X=35655 $Y=30285
X5796 355 346 VDD 373 376 VSS 344 670 AOI221_X1 $T=35960 20600 1 0 $X=35845 $Y=19085
X5797 351 324 VDD 371 387 VSS 514 918 AOI221_X1 $T=36530 34600 1 0 $X=36415 $Y=33085
X5798 394 346 VDD 373 390 VSS 344 393 AOI221_X1 $T=38240 20600 0 180 $X=36985 $Y=19085
X5799 670 821 VDD 403 408 VSS 920 421 AOI221_X1 $T=38810 20600 0 0 $X=38695 $Y=20485
X5800 420 461 VDD 434 429 VSS 889 sum[5] AOI221_X1 $T=42230 45800 1 0 $X=42115 $Y=44285
X5801 429 837 VDD 444 420 VSS 889 sum[6] AOI221_X1 $T=44320 45800 1 180 $X=43065 $Y=45685
X5802 420 837 VDD 456 459 VSS 429 sum[7] AOI221_X1 $T=44320 45800 0 0 $X=44205 $Y=45685
X5803 420 836 VDD 478 429 VSS 453 sum[19] AOI221_X1 $T=46790 20600 1 180 $X=45535 $Y=20485
X5804 420 712 VDD 470 429 VSS 836 sum[18] AOI221_X1 $T=45650 23400 1 0 $X=45535 $Y=21885
X5805 429 712 VDD 471 479 VSS 420 sum[17] AOI221_X1 $T=45650 23400 0 0 $X=45535 $Y=23285
X5806 420 706 VDD 472 429 VSS 846 sum[15] AOI221_X1 $T=45650 26200 0 0 $X=45535 $Y=26085
X5807 487 429 VDD 473 420 VSS 533 sum[13] AOI221_X1 $T=45650 31800 1 0 $X=45535 $Y=30285
X5808 420 488 VDD 474 429 VSS 717 sum[11] AOI221_X1 $T=45650 37400 1 0 $X=45535 $Y=35885
X5809 420 467 VDD 475 480 VSS 429 sum[9] AOI221_X1 $T=45650 40200 0 0 $X=45535 $Y=40085
X5810 420 459 VDD 476 467 VSS 429 sum[8] AOI221_X1 $T=45650 45800 1 0 $X=45535 $Y=44285
X5811 429 706 VDD 482 487 VSS 420 sum[14] AOI221_X1 $T=46030 29000 0 0 $X=45915 $Y=28885
X5812 420 717 VDD 483 429 VSS 533 sum[12] AOI221_X1 $T=46030 34600 1 0 $X=45915 $Y=33085
X5813 420 480 VDD 484 488 VSS 429 sum[10] AOI221_X1 $T=46030 40200 1 0 $X=45915 $Y=38685
X5814 372 402 VSS 396 398 VDD 401 sum[2] OAI221_X1 $T=37670 37400 0 0 $X=37555 $Y=37285
X5815 714 401 VSS 443 446 VDD 398 sum[3] OAI221_X1 $T=43370 37400 1 0 $X=43255 $Y=35885
X5816 714 453 VSS 452 398 VDD 481 sum[20] OAI221_X1 $T=44890 20600 0 180 $X=43635 $Y=19085
X5817 714 446 VSS 458 461 VDD 398 sum[4] OAI221_X1 $T=44510 37400 1 0 $X=44395 $Y=35885
X5818 714 846 VSS 486 398 VDD 479 sum[16] OAI221_X1 $T=47170 26200 0 180 $X=45915 $Y=24685
X5819 42 36 51 45 VSS VDD VSS OAI21_X1 $T=3090 45800 0 0 $X=2975 $Y=45685
X5820 537 54 539 64 VSS VDD VSS OAI21_X1 $T=4990 6600 0 0 $X=4875 $Y=6485
X5821 68 65 55 544 VSS VDD VSS OAI21_X1 $T=5750 17800 0 0 $X=5635 $Y=17685
X5822 53 56 63 86 VSS VDD VSS OAI21_X1 $T=6510 34600 0 180 $X=5635 $Y=33085
X5823 76 66 91 80 VSS VDD VSS OAI21_X1 $T=5750 43000 1 0 $X=5635 $Y=41485
X5824 537 71 732 499 VSS VDD VSS OAI21_X1 $T=7080 9400 1 180 $X=6205 $Y=9285
X5825 497 105 856 117 VSS VDD VSS OAI21_X1 $T=8600 9400 1 0 $X=8485 $Y=7885
X5826 574 109 499 117 VSS VDD VSS OAI21_X1 $T=9360 9400 1 0 $X=9245 $Y=7885
X5827 132 136 141 135 VSS VDD VSS OAI21_X1 $T=11070 40200 1 0 $X=10955 $Y=38685
X5828 148 150 160 173 VSS VDD VSS OAI21_X1 $T=14490 34600 0 180 $X=13615 $Y=33085
X5829 b[23] b[24] 151 b[25] VSS VDD VSS OAI21_X1 $T=13920 3800 0 0 $X=13805 $Y=3685
X5830 108 159 580 505 VSS VDD VSS OAI21_X1 $T=14870 20600 1 180 $X=13995 $Y=20485
X5831 74 140 179 569 VSS VDD VSS OAI21_X1 $T=15060 9400 1 180 $X=14185 $Y=9285
X5832 74 140 175 574 VSS VDD VSS OAI21_X1 $T=15060 9400 0 0 $X=14945 $Y=9285
X5833 166 174 177 170 VSS VDD VSS OAI21_X1 $T=15630 40200 1 0 $X=15515 $Y=38685
X5834 232 236 245 227 VSS VDD VSS OAI21_X1 $T=22660 12200 0 180 $X=21785 $Y=10685
X5835 265 272 278 267 VSS VDD VSS OAI21_X1 $T=25510 45800 1 0 $X=25395 $Y=44285
X5836 257 255 281 342 VSS VDD VSS OAI21_X1 $T=26650 37400 1 180 $X=25775 $Y=37285
X5837 312 311 952 313 VSS VDD VSS OAI21_X1 $T=29310 15000 0 0 $X=29195 $Y=14885
X5838 298 321 326 297 VSS VDD VSS OAI21_X1 $T=30830 45800 0 180 $X=29955 $Y=44285
X5839 901 332 874 938 VSS VDD VSS OAI21_X1 $T=31780 31800 1 180 $X=30905 $Y=31685
X5840 516 337 sum[31] 799 VSS VDD VSS OAI21_X1 $T=31970 3800 1 0 $X=31855 $Y=2285
X5841 341 339 389 650 VSS VDD VSS OAI21_X1 $T=33300 17800 1 180 $X=32425 $Y=17685
X5842 878 343 903 649 VSS VDD VSS OAI21_X1 $T=33490 43000 0 180 $X=32615 $Y=41485
X5843 385 308 692 906 VSS VDD VSS OAI21_X1 $T=34060 34600 0 0 $X=33945 $Y=34485
X5844 656 357 676 661 VSS VDD VSS OAI21_X1 $T=34440 20600 0 0 $X=34325 $Y=20485
X5845 524 363 660 347 VSS VDD VSS OAI21_X1 $T=34820 34600 0 0 $X=34705 $Y=34485
X5846 941 388 907 672 VSS VDD 975 OAI21_X1 $T=36910 1000 0 0 $X=36795 $Y=885
X5847 383 386 sum[1] 671 VSS VDD VSS OAI21_X1 $T=37670 37400 1 180 $X=36795 $Y=37285
X5848 679 387 688 817 VSS VDD VSS OAI21_X1 $T=38430 34600 0 180 $X=37555 $Y=33085
X5849 400 397 435 676 VSS VDD VSS OAI21_X1 $T=37860 17800 0 0 $X=37745 $Y=17685
X5850 884 399 819 527 VSS VDD VSS OAI21_X1 $T=37860 43000 0 0 $X=37745 $Y=42885
X5851 912 335 400 911 VSS VDD VSS OAI21_X1 $T=39000 12200 1 180 $X=38125 $Y=12085
X5852 385 334 678 528 VSS VDD VSS OAI21_X1 $T=38240 29000 1 0 $X=38125 $Y=27485
X5853 679 257 427 681 VSS VDD VSS OAI21_X1 $T=38810 31800 0 0 $X=38695 $Y=31685
X5854 689 426 442 687 VSS VDD VSS OAI21_X1 $T=41090 26200 1 0 $X=40975 $Y=24685
X5855 419 427 827 829 VSS VDD VSS OAI21_X1 $T=41090 31800 1 0 $X=40975 $Y=30285
X5856 419 436 922 697 VSS VDD VSS OAI21_X1 $T=42420 31800 0 0 $X=42305 $Y=31685
X5857 371 436 835 699 VSS VDD VSS OAI21_X1 $T=43180 34600 0 0 $X=43065 $Y=34485
X5858 530 442 453 950 VSS VDD VSS OAI21_X1 $T=44320 20600 1 180 $X=43445 $Y=20485
X5859 530 445 479 704 VSS VDD VSS OAI21_X1 $T=44510 26200 1 180 $X=43635 $Y=26085
X5860 408 448 837 708 VSS VDD VSS OAI21_X1 $T=43750 43000 0 0 $X=43635 $Y=42885
X5861 530 462 712 944 VSS VDD VSS OAI21_X1 $T=44890 23400 0 0 $X=44775 $Y=23285
X5862 408 468 459 715 VSS VDD VSS OAI21_X1 $T=45460 43000 0 0 $X=45345 $Y=42885
X5863 714 481 sum[21] 721 VSS VDD VSS OAI21_X1 $T=46030 17800 0 0 $X=45915 $Y=17685
X6025 125 122 VDD 489 554 541 VSS AOI22_X1 $T=4800 17800 0 0 $X=4685 $Y=17685
X6026 59 121 VDD 540 61 541 VSS AOI22_X1 $T=5940 17800 0 180 $X=4875 $Y=16285
X6027 119 122 VDD 726 854 541 VSS AOI22_X1 $T=4990 23400 1 0 $X=4875 $Y=21885
X6028 727 122 VDD 923 93 541 VSS AOI22_X1 $T=4990 26200 1 0 $X=4875 $Y=24685
X6029 115 551 VDD 81 729 52 VSS AOI22_X1 $T=4990 26200 0 0 $X=4875 $Y=26085
X6030 129 551 VDD 725 733 111 VSS AOI22_X1 $T=7080 12200 0 0 $X=6965 $Y=12085
X6031 68 730 VDD 552 925 111 VSS AOI22_X1 $T=7080 29000 1 0 $X=6965 $Y=27485
X6032 925 549 VDD 137 859 74 VSS AOI22_X1 $T=7460 26200 0 0 $X=7345 $Y=26085
X6033 504 560 VDD 567 753 563 VSS AOI22_X1 $T=12780 15000 0 0 $X=12665 $Y=14885
X6034 111 748 VDD 559 566 85 VSS AOI22_X1 $T=12780 17800 1 0 $X=12665 $Y=16285
X6035 504 567 VDD 140 929 565 VSS AOI22_X1 $T=13920 12200 1 180 $X=12855 $Y=12085
X6036 563 560 VDD 159 572 108 VSS AOI22_X1 $T=12970 17800 0 0 $X=12855 $Y=17685
X6037 110 565 VDD 567 576 133 VSS AOI22_X1 $T=14110 15000 0 180 $X=13045 $Y=13485
X6038 926 756 VDD 573 583 582 VSS AOI22_X1 $T=16200 45800 0 0 $X=16085 $Y=45685
X6039 898 774 VDD 599 606 604 VSS AOI22_X1 $T=22280 31800 0 0 $X=22165 $Y=31685
X6040 608 775 VDD 934 953 782 VSS AOI22_X1 $T=24560 20600 1 0 $X=24445 $Y=19085
X6041 637 598 VDD 509 802 793 VSS AOI22_X1 $T=31020 9400 1 0 $X=30905 $Y=7885
X6042 631 344 VDD 312 807 346 VSS AOI22_X1 $T=31970 20600 1 0 $X=31855 $Y=19085
X6043 257 514 VDD 299 651 346 VSS AOI22_X1 $T=32540 29000 1 0 $X=32425 $Y=27485
X6044 632 344 VDD 314 905 346 VSS AOI22_X1 $T=32920 23400 0 0 $X=32805 $Y=23285
X6045 514 654 VDD 308 879 351 VSS AOI22_X1 $T=33110 34600 1 0 $X=32995 $Y=33085
X6046 514 698 VDD 325 658 351 VSS AOI22_X1 $T=34060 34600 1 0 $X=33945 $Y=33085
X6047 796 808 VDD 804 664 663 VSS AOI22_X1 $T=34440 6600 0 0 $X=34325 $Y=6485
X6048 428 271 VDD 698 396 667 VSS AOI22_X1 $T=35010 37400 0 0 $X=34895 $Y=37285
X6049 314 428 VDD 299 486 424 VSS AOI22_X1 $T=35770 23400 0 0 $X=35655 $Y=23285
X6050 257 667 VDD 342 671 428 VSS AOI22_X1 $T=36910 37400 1 180 $X=35845 $Y=37285
X6051 514 381 VDD 322 821 351 VSS AOI22_X1 $T=37290 29000 0 180 $X=36225 $Y=27485
X6052 514 815 VDD 334 395 351 VSS AOI22_X1 $T=37290 29000 1 0 $X=37175 $Y=27485
X6053 428 290 VDD 387 443 424 VSS AOI22_X1 $T=38810 37400 0 0 $X=38695 $Y=37285
X6054 428 298 VDD 374 458 424 VSS AOI22_X1 $T=39760 37400 0 0 $X=39645 $Y=37285
X6055 694 387 VDD 515 710 377 VSS AOI22_X1 $T=40520 40200 0 0 $X=40405 $Y=40085
X6056 355 428 VDD 340 452 424 VSS AOI22_X1 $T=40900 15000 1 0 $X=40785 $Y=13485
X6057 257 694 VDD 374 826 377 VSS AOI22_X1 $T=41850 40200 0 180 $X=40785 $Y=38685
X6058 257 433 VDD 654 401 412 VSS AOI22_X1 $T=41470 37400 1 0 $X=41355 $Y=35885
X6059 694 698 VDD 381 701 377 VSS AOI22_X1 $T=41470 40200 0 0 $X=41355 $Y=40085
X6060 654 433 VDD 530 461 833 VSS AOI22_X1 $T=42230 40200 1 0 $X=42115 $Y=38685
X6061 433 698 VDD 387 446 412 VSS AOI22_X1 $T=42420 37400 1 0 $X=42305 $Y=35885
X6062 694 654 VDD 815 707 377 VSS AOI22_X1 $T=42420 40200 0 0 $X=42305 $Y=40085
X6063 696 831 VDD 419 440 703 VSS AOI22_X1 $T=42800 26200 0 0 $X=42685 $Y=26085
X6064 530 445 VDD 705 706 827 VSS AOI22_X1 $T=44510 29000 0 180 $X=43445 $Y=27485
X6065 922 705 VDD 530 846 462 VSS AOI22_X1 $T=44510 29000 1 0 $X=44395 $Y=27485
X6066 705 682 VDD 922 487 466 VSS AOI22_X1 $T=45650 31800 1 180 $X=44585 $Y=31685
X6067 448 408 VDD 825 467 466 VSS AOI22_X1 $T=44700 40200 0 0 $X=44585 $Y=40085
X6068 466 460 VDD 825 488 705 VSS AOI22_X1 $T=44890 34600 0 0 $X=44775 $Y=34485
X6069 468 408 VDD 835 480 466 VSS AOI22_X1 $T=45080 40200 1 0 $X=44965 $Y=38685
X6070 705 835 VDD 466 717 682 VSS AOI22_X1 $T=45840 34600 0 0 $X=45725 $Y=34485
X6071 b[16] 18 a[16] VSS VDD 79 VSS MUX2_X1 $T=2330 17800 1 180 $X=885 $Y=17685
X6072 a[5] 37 b[5] VSS VDD 42 VSS MUX2_X1 $T=2330 23400 0 180 $X=885 $Y=21885
X6073 a[4] 37 b[4] VSS VDD 44 VSS MUX2_X1 $T=2330 26200 1 180 $X=885 $Y=26085
X6074 a[3] 37 b[3] VSS VDD 57 VSS MUX2_X1 $T=2330 31800 1 180 $X=885 $Y=31685
X6075 a[10] 37 b[10] VSS VDD 99 VSS MUX2_X1 $T=1000 37400 1 0 $X=885 $Y=35885
X6076 b[6] 18 a[6] VSS VDD 489 VSS MUX2_X1 $T=2330 40200 1 180 $X=885 $Y=40085
X6077 a[15] 37 b[15] VSS VDD 205 VSS MUX2_X1 $T=3660 15000 1 180 $X=2215 $Y=14885
X6078 a[14] 37 b[14] VSS VDD 214 VSS MUX2_X1 $T=3660 17800 0 180 $X=2215 $Y=16285
X6079 b[14] 18 a[14] VSS VDD 125 VSS MUX2_X1 $T=2330 17800 0 0 $X=2215 $Y=17685
X6080 a[16] 37 b[16] VSS VDD 184 VSS MUX2_X1 $T=3660 20600 0 180 $X=2215 $Y=19085
X6081 b[11] 18 a[11] VSS VDD 49 VSS MUX2_X1 $T=3660 29000 0 180 $X=2215 $Y=27485
X6082 b[3] 18 a[3] VSS VDD VDD VSS MUX2_X1 $T=3660 31800 0 180 $X=2215 $Y=30285
X6083 b[1] 18 a[1] VSS VDD 62 VSS MUX2_X1 $T=3660 31800 1 180 $X=2215 $Y=31685
X6084 b[9] 18 a[9] VSS VDD 81 VSS MUX2_X1 $T=3660 37400 0 180 $X=2215 $Y=35885
X6085 b[7] 18 a[7] VSS VDD 535 VSS MUX2_X1 $T=3660 40200 0 180 $X=2215 $Y=38685
X6086 b[8] 18 a[8] VSS VDD 102 VSS MUX2_X1 $T=3660 40200 1 180 $X=2215 $Y=40085
X6087 49 68 43 VSS VDD 94 VSS MUX2_X1 $T=4990 15000 0 180 $X=3545 $Y=13485
X6088 a[17] 37 b[17] VSS VDD 189 VSS MUX2_X1 $T=3660 20600 1 0 $X=3545 $Y=19085
X6089 b[0] 18 a[0] VSS VDD 552 VSS MUX2_X1 $T=4990 31800 0 180 $X=3545 $Y=30285
X6090 a[0] 37 b[0] VSS VDD 53 VSS MUX2_X1 $T=3660 31800 0 0 $X=3545 $Y=31685
X6091 70 638 42 VSS VDD 914 VSS MUX2_X1 $T=6700 45800 1 180 $X=5255 $Y=45685
X6092 73 638 44 VSS VDD 924 VSS MUX2_X1 $T=6890 40200 0 180 $X=5445 $Y=38685
X6093 75 638 86 VSS VDD 897 VSS MUX2_X1 $T=6510 34600 0 0 $X=6395 $Y=34485
X6094 82 74 89 VSS VDD 927 VSS MUX2_X1 $T=6890 29000 0 0 $X=6775 $Y=28885
X6095 90 638 99 VSS VDD 734 VSS MUX2_X1 $T=7460 40200 1 0 $X=7345 $Y=38685
X6096 92 638 80 VSS VDD 735 VSS MUX2_X1 $T=7460 43000 1 0 $X=7345 $Y=41485
X6097 96 638 103 VSS VDD 898 VSS MUX2_X1 $T=7840 31800 0 0 $X=7725 $Y=31685
X6098 100 638 45 VSS VDD 736 VSS MUX2_X1 $T=8030 45800 0 0 $X=7915 $Y=45685
X6099 107 108 89 VSS VDD 745 VSS MUX2_X1 $T=9550 29000 1 180 $X=8105 $Y=28885
X6100 a[30] 18 b[30] VSS VDD 737 975 MUX2_X1 $T=10880 1000 1 180 $X=9435 $Y=885
X6101 112 108 107 VSS VDD 127 VSS MUX2_X1 $T=9550 29000 0 0 $X=9435 $Y=28885
X6102 116 139 123 VSS VDD 142 VSS MUX2_X1 $T=9740 37400 0 0 $X=9625 $Y=37285
X6103 134 108 126 VSS VDD 500 VSS MUX2_X1 $T=11640 26200 1 180 $X=10195 $Y=26085
X6104 129 68 118 VSS VDD 133 VSS MUX2_X1 $T=10690 15000 1 0 $X=10575 $Y=13485
X6105 137 74 126 VSS VDD 742 VSS MUX2_X1 $T=12020 29000 0 180 $X=10575 $Y=27485
X6106 138 139 132 VSS VDD 739 VSS MUX2_X1 $T=12020 40200 1 180 $X=10575 $Y=40085
X6107 131 638 56 VSS VDD 746 VSS MUX2_X1 $T=10880 34600 0 0 $X=10765 $Y=34485
X6108 115 68 140 VSS VDD 563 VSS MUX2_X1 $T=11260 20600 0 0 $X=11145 $Y=20485
X6109 79 74 129 VSS VDD 748 VSS MUX2_X1 $T=11450 17800 1 0 $X=11335 $Y=16285
X6110 79 68 110 VSS VDD 155 VSS MUX2_X1 $T=11450 20600 1 0 $X=11335 $Y=19085
X6111 145 108 134 VSS VDD 749 VSS MUX2_X1 $T=12970 26200 1 180 $X=11525 $Y=26085
X6112 147 108 112 VSS VDD 928 VSS MUX2_X1 $T=13350 29000 0 180 $X=11905 $Y=27485
X6113 144 139 135 VSS VDD 747 VSS MUX2_X1 $T=12020 40200 0 0 $X=11905 $Y=40085
X6114 154 108 145 VSS VDD 570 VSS MUX2_X1 $T=14300 26200 1 180 $X=12855 $Y=26085
X6115 152 74 156 VSS VDD 751 VSS MUX2_X1 $T=13350 23400 0 0 $X=13235 $Y=23285
X6116 152 108 147 VSS VDD 752 VSS MUX2_X1 $T=13350 29000 1 0 $X=13235 $Y=27485
X6117 154 74 163 VSS VDD 754 VSS MUX2_X1 $T=14300 26200 1 0 $X=14185 $Y=24685
X6118 162 108 163 VSS VDD 930 VSS MUX2_X1 $T=14870 23400 1 0 $X=14755 $Y=21885
X6119 165 139 173 VSS VDD 767 VSS MUX2_X1 $T=15250 34600 0 0 $X=15135 $Y=34485
X6120 167 139 166 VSS VDD 188 VSS MUX2_X1 $T=15250 43000 0 0 $X=15135 $Y=42885
X6121 171 139 157 VSS VDD 756 VSS MUX2_X1 $T=15440 43000 1 0 $X=15325 $Y=41485
X6122 a[24] 18 b[24] VSS VDD 439 VSS MUX2_X1 $T=17150 6600 0 180 $X=15705 $Y=5085
X6123 a[25] 18 b[25] VSS VDD 463 VSS MUX2_X1 $T=18100 3800 1 180 $X=16655 $Y=3685
X6124 181 139 150 VSS VDD 757 VSS MUX2_X1 $T=16770 34600 1 0 $X=16655 $Y=33085
X6125 183 139 170 VSS VDD 931 VSS MUX2_X1 $T=17150 40200 1 0 $X=17035 $Y=38685
X6126 a[28] 18 b[28] VSS VDD 413 975 MUX2_X1 $T=18670 1000 1 180 $X=17225 $Y=885
X6127 197 638 189 VSS VDD 899 VSS MUX2_X1 $T=19050 15000 1 180 $X=17605 $Y=14885
X6128 b[19] 18 a[19] VSS VDD 60 VSS MUX2_X1 $T=19240 3800 0 180 $X=17795 $Y=2285
X6129 194 139 202 VSS VDD 765 VSS MUX2_X1 $T=18100 37400 0 0 $X=17985 $Y=37285
X6130 200 638 205 VSS VDD 608 VSS MUX2_X1 $T=18670 20600 0 0 $X=18555 $Y=20485
X6131 215 139 208 VSS VDD 808 VSS MUX2_X1 $T=20570 6600 1 180 $X=19125 $Y=6485
X6132 209 638 184 VSS VDD 613 VSS MUX2_X1 $T=19430 17800 0 0 $X=19315 $Y=17685
X6133 211 638 196 VSS VDD 779 VSS MUX2_X1 $T=19620 12200 1 0 $X=19505 $Y=10685
X6134 217 139 225 VSS VDD 598 VSS MUX2_X1 $T=20570 6600 0 0 $X=20455 $Y=6485
X6135 221 139 230 VSS VDD 774 VSS MUX2_X1 $T=20570 31800 1 0 $X=20455 $Y=30285
X6136 a[29] 18 b[29] VSS VDD 932 975 MUX2_X1 $T=23040 1000 1 180 $X=21595 $Y=885
X6137 238 139 246 VSS VDD 775 VSS MUX2_X1 $T=22090 20600 1 0 $X=21975 $Y=19085
X6138 249 139 227 VSS VDD 935 VSS MUX2_X1 $T=23420 12200 1 0 $X=23305 $Y=10685
X6139 a[22] 37 b[22] VSS VDD 317 VSS MUX2_X1 $T=23610 3800 1 0 $X=23495 $Y=2285
X6140 263 638 260 VSS VDD 626 VSS MUX2_X1 $T=25890 6600 1 180 $X=24445 $Y=6485
X6141 264 139 273 VSS VDD 937 VSS MUX2_X1 $T=25320 9400 1 0 $X=25205 $Y=7885
X6142 266 139 276 VSS VDD 292 VSS MUX2_X1 $T=25510 9400 0 0 $X=25395 $Y=9285
X6143 279 638 283 VSS VDD 788 VSS MUX2_X1 $T=26460 6600 0 0 $X=26345 $Y=6485
X6144 a[20] 37 b[20] VSS VDD 260 VSS MUX2_X1 $T=26840 3800 1 0 $X=26725 $Y=2285
X6145 293 333 288 VSS VDD 308 VSS MUX2_X1 $T=28550 40200 1 180 $X=27105 $Y=40085
X6146 269 333 289 VSS VDD 324 VSS MUX2_X1 $T=28740 37400 0 180 $X=27295 $Y=35885
X6147 b[20] 18 a[20] VSS VDD 110 975 MUX2_X1 $T=28930 1000 1 180 $X=27485 $Y=885
X6148 265 333 301 VSS VDD 336 VSS MUX2_X1 $T=28170 45800 0 0 $X=28055 $Y=45685
X6149 267 333 306 VSS VDD 325 VSS MUX2_X1 $T=28550 43000 0 0 $X=28435 $Y=42885
X6150 255 333 302 VSS VDD 698 VSS MUX2_X1 $T=30070 34600 0 180 $X=28625 $Y=33085
X6151 269 318 308 VSS VDD 634 VSS MUX2_X1 $T=28740 37400 1 0 $X=28625 $Y=35885
X6152 305 333 315 VSS VDD 334 VSS MUX2_X1 $T=29120 29000 1 0 $X=29005 $Y=27485
X6153 290 333 316 VSS VDD 374 VSS MUX2_X1 $T=29120 40200 1 0 $X=29005 $Y=38685
X6154 307 638 317 VSS VDD 637 VSS MUX2_X1 $T=29310 6600 1 0 $X=29195 $Y=5085
X6155 274 318 324 VSS VDD 332 VSS MUX2_X1 $T=30070 34600 1 0 $X=29955 $Y=33085
X6156 293 318 325 VSS VDD 643 VSS MUX2_X1 $T=30070 40200 0 0 $X=29955 $Y=40085
X6157 328 318 334 VSS VDD 511 VSS MUX2_X1 $T=30830 26200 0 0 $X=30715 $Y=26085
X6158 267 318 336 VSS VDD 513 VSS MUX2_X1 $T=31400 43000 1 0 $X=31285 $Y=41485
X6159 342 348 338 VSS VDD 654 VSS MUX2_X1 $T=33300 40200 0 180 $X=31855 $Y=38685
X6160 275 348 794 VSS VDD 515 VSS MUX2_X1 $T=34060 45800 1 180 $X=32615 $Y=45685
X6161 298 348 352 VSS VDD 381 VSS MUX2_X1 $T=33110 43000 0 0 $X=32995 $Y=42885
X6162 354 388 360 VSS VDD sum[29] VSS MUX2_X1 $T=34250 3800 1 0 $X=34135 $Y=2285
X6163 297 348 384 VSS VDD 815 VSS MUX2_X1 $T=36150 45800 0 0 $X=36035 $Y=45685
X6164 322 385 381 VSS VDD 830 VSS MUX2_X1 $T=37670 29000 1 180 $X=36225 $Y=28885
X6165 297 318 381 VSS VDD 378 VSS MUX2_X1 $T=38050 45800 1 0 $X=37935 $Y=44285
X6166 290 318 387 VSS VDD 399 VSS MUX2_X1 $T=40330 43000 0 180 $X=38885 $Y=41485
X6167 405 388 410 VSS VDD sum[28] VSS MUX2_X1 $T=39190 3800 1 0 $X=39075 $Y=2285
X6168 a[26] 18 b[26] VSS VDD 465 VSS MUX2_X1 $T=41850 3800 0 180 $X=40405 $Y=2285
X6169 418 388 423 VSS VDD sum[23] VSS MUX2_X1 $T=40520 12200 1 0 $X=40405 $Y=10685
X6170 a[27] 18 b[27] VSS VDD 709 975 MUX2_X1 $T=41090 1000 0 0 $X=40975 $Y=885
X6171 431 530 437 VSS VDD 481 VSS MUX2_X1 $T=42230 20600 0 0 $X=42115 $Y=20485
X6172 431 408 440 VSS VDD 836 VSS MUX2_X1 $T=42800 23400 1 0 $X=42685 $Y=21885
X6173 447 388 454 VSS VDD sum[27] 975 MUX2_X1 $T=43940 1000 0 0 $X=43825 $Y=885
X6174 469 388 485 VSS VDD sum[24] VSS MUX2_X1 $T=45840 12200 1 0 $X=45725 $Y=10685
X6183 VSS 849 893 35 VDD VSS XNOR2_X1 $T=2900 9400 1 0 $X=2785 $Y=7885
X6184 VSS 543 728 64 VDD VSS XNOR2_X1 $T=6700 9400 0 180 $X=5445 $Y=7885
X6185 VSS 103 96 83 VDD VSS XNOR2_X1 $T=6700 31800 0 0 $X=6585 $Y=31685
X6186 VSS b[30] 851 104 VDD 975 XNOR2_X1 $T=9550 1000 1 180 $X=8295 $Y=885
X6187 VSS 205 200 186 VDD VSS XNOR2_X1 $T=17530 20600 0 0 $X=17415 $Y=20485
X6188 VSS 214 206 190 VDD VSS XNOR2_X1 $T=17720 23400 0 0 $X=17605 $Y=23285
X6189 VSS 208 215 195 VDD VSS XNOR2_X1 $T=18100 6600 0 0 $X=17985 $Y=6485
X6190 VSS 196 211 896 VDD VSS XNOR2_X1 $T=18480 12200 1 0 $X=18365 $Y=10685
X6191 VSS 230 221 213 VDD VSS XNOR2_X1 $T=19430 31800 1 0 $X=19315 $Y=30285
X6192 VSS 247 239 223 VDD VSS XNOR2_X1 $T=20760 3800 0 0 $X=20645 $Y=3685
X6193 VSS 225 217 226 VDD VSS XNOR2_X1 $T=21900 9400 1 180 $X=20645 $Y=9285
X6194 VSS 246 238 863 VDD VSS XNOR2_X1 $T=20760 20600 0 0 $X=20645 $Y=20485
X6195 VSS 164 219 228 VDD VSS XNOR2_X1 $T=21900 23400 1 180 $X=20645 $Y=23285
X6196 VSS 273 264 243 VDD VSS XNOR2_X1 $T=22280 9400 1 0 $X=22165 $Y=7885
X6197 VSS 269 289 270 VDD VSS XNOR2_X1 $T=25700 34600 0 0 $X=25585 $Y=34485
X6198 VSS 305 315 285 VDD VSS XNOR2_X1 $T=26840 26200 0 0 $X=26725 $Y=26085
X6199 VSS 317 307 294 VDD VSS XNOR2_X1 $T=27980 3800 0 0 $X=27865 $Y=3685
X6200 VSS 328 792 304 VDD VSS XNOR2_X1 $T=28930 26200 1 0 $X=28815 $Y=24685
X6201 VSS 737 sum[30] 907 VDD 975 XNOR2_X1 $T=33870 1000 0 0 $X=33755 $Y=885
X6202 VSS 516 335 366 VDD VSS XNOR2_X1 $T=36150 12200 1 180 $X=34895 $Y=12085
X6203 VSS 355 376 369 VDD VSS XNOR2_X1 $T=36530 12200 0 180 $X=35275 $Y=10685
X6204 VSS 803 673 379 VDD VSS XNOR2_X1 $T=36340 3800 0 0 $X=36225 $Y=3685
X6205 VSS 409 675 407 VDD VSS XNOR2_X1 $T=39950 9400 1 180 $X=38695 $Y=9285
X6206 VSS 394 390 411 VDD VSS XNOR2_X1 $T=40520 12200 0 180 $X=39265 $Y=10685
X6207 VSS 371 891 432 VDD VSS XNOR2_X1 $T=42230 17800 1 0 $X=42115 $Y=16285
X6208 VSS 523 890 441 VDD VSS XNOR2_X1 $T=44320 15000 0 180 $X=43065 $Y=13485
X6209 VSS 530 892 435 VDD VSS XNOR2_X1 $T=45650 15000 1 0 $X=45535 $Y=13485
X6958 VSS VDD a[23] 18 b[23] 690 ICV_14 $T=16580 6600 0 0 $X=16465 $Y=6485
X6959 VSS VDD 187 638 176 602 ICV_14 $T=17530 29000 0 0 $X=17415 $Y=28885
X6960 VSS VDD 271 333 319 387 ICV_14 $T=29120 37400 0 0 $X=29005 $Y=37285
X6961 VSS VDD 255 318 257 816 ICV_14 $T=29310 34600 0 0 $X=29195 $Y=34485
X6962 VSS VDD 305 318 322 642 ICV_14 $T=29690 29000 0 0 $X=29575 $Y=28885
X6963 VSS VDD 340 333 345 657 ICV_14 $T=32540 15000 0 0 $X=32425 $Y=14885
X6964 VSS VDD 449 388 457 sum[26] ICV_14 $T=43940 6600 1 0 $X=43825 $Y=5085
X6965 VSS VDD 464 388 477 sum[25] ICV_14 $T=45270 9400 0 0 $X=45155 $Y=9285
X6966 574 a[23] b[23] VSS VDD 130 VSS HA_X1 $T=14490 9400 0 180 $X=12475 $Y=7885
X6967 354 666 932 VSS VDD 941 975 HA_X1 $T=35010 1000 0 0 $X=34895 $Y=885
X6968 405 724 413 VSS VDD 666 975 HA_X1 $T=39190 1000 0 0 $X=39075 $Y=885
X6969 418 690 428 VSS VDD 700 VSS HA_X1 $T=39950 9400 0 0 $X=39835 $Y=9285
X6970 423 690 435 VSS VDD 451 VSS HA_X1 $T=41850 12200 0 0 $X=41735 $Y=12085
X6971 469 700 439 VSS VDD 529 VSS HA_X1 $T=42230 9400 0 0 $X=42115 $Y=9285
X6972 449 711 465 VSS VDD 713 VSS HA_X1 $T=44890 3800 0 0 $X=44775 $Y=3685
X6973 464 529 463 VSS VDD 711 VSS HA_X1 $T=46790 6600 1 180 $X=44775 $Y=6485
X6974 447 713 709 VSS VDD 724 975 HA_X1 $T=45270 1000 0 0 $X=45155 $Y=885
X7000 59 94 498 VDD 101 152 VSS OAI211_X1 $T=7650 15000 1 0 $X=7535 $Y=13485
X7001 68 121 955 VDD 128 159 VSS OAI211_X1 $T=10120 17800 1 0 $X=10005 $Y=16285
X7002 417 414 686 VDD 948 823 VSS OAI211_X1 $T=40710 23400 0 180 $X=39645 $Y=21885
X7003 530 460 691 VDD 455 533 VSS OAI211_X1 $T=45650 31800 0 180 $X=44585 $Y=30285
X7045 537 VSS VDD 492 INV_X1 $T=1760 9400 1 0 $X=1645 $Y=7885
X7046 535 VSS VDD 540 INV_X1 $T=4420 29000 0 0 $X=4305 $Y=28885
X7047 543 VSS VDD 54 INV_X1 $T=6130 6600 1 180 $X=5635 $Y=6485
X7048 545 VSS VDD 498 INV_X1 $T=6130 15000 0 180 $X=5635 $Y=13485
X7049 729 VSS VDD 69 INV_X1 $T=5940 26200 0 0 $X=5825 $Y=26085
X7050 497 VSS VDD 71 INV_X1 $T=7080 9400 0 180 $X=6585 $Y=7885
X7051 122 VSS VDD 548 INV_X1 $T=6700 23400 1 0 $X=6585 $Y=21885
X7052 103 VSS VDD 949 INV_X1 $T=6890 31800 1 0 $X=6775 $Y=30285
X7053 68 VSS VDD 87 INV_X1 $T=7460 15000 0 0 $X=7345 $Y=14885
X7054 733 VSS VDD 95 INV_X1 $T=8600 15000 1 0 $X=8485 $Y=13485
X7055 556 VSS VDD 504 INV_X1 $T=10690 12200 0 0 $X=10575 $Y=12085
X7056 859 VSS VDD 740 INV_X1 $T=10880 29000 0 0 $X=10765 $Y=28885
X7057 52 VSS VDD 955 INV_X1 $T=11450 17800 0 180 $X=10955 $Y=16285
X7058 744 VSS VDD 564 INV_X1 $T=11830 45800 1 0 $X=11715 $Y=44285
X7059 574 VSS VDD 569 INV_X1 $T=13350 9400 1 180 $X=12855 $Y=9285
X7060 568 VSS VDD 582 INV_X1 $T=14110 45800 0 0 $X=13995 $Y=45685
X7061 74 VSS VDD 108 INV_X1 $T=15060 15000 0 0 $X=14945 $Y=14885
X7062 205 VSS VDD 579 INV_X1 $T=16390 17800 0 0 $X=16275 $Y=17685
X7063 583 VSS VDD 204 INV_X1 $T=17150 45800 0 0 $X=17035 $Y=45685
X7064 246 VSS VDD 763 INV_X1 $T=19430 20600 1 0 $X=19315 $Y=19085
X7065 590 VSS VDD 770 INV_X1 $T=19430 40200 0 0 $X=19315 $Y=40085
X7066 230 VSS VDD 862 INV_X1 $T=20000 29000 1 180 $X=19505 $Y=28885
X7067 865 VSS VDD 771 INV_X1 $T=20570 34600 0 0 $X=20455 $Y=34485
X7068 222 VSS VDD 595 INV_X1 $T=20760 37400 1 0 $X=20645 $Y=35885
X7069 866 VSS VDD 772 INV_X1 $T=21140 40200 1 180 $X=20645 $Y=40085
X7070 247 VSS VDD 597 INV_X1 $T=21520 6600 1 0 $X=21405 $Y=5085
X7071 596 VSS VDD 604 INV_X1 $T=21520 37400 0 0 $X=21405 $Y=37285
X7072 606 VSS VDD 256 INV_X1 $T=23420 31800 0 0 $X=23305 $Y=31685
X7073 867 VSS VDD 617 INV_X1 $T=23990 26200 0 0 $X=23875 $Y=26085
X7074 869 VSS VDD 782 INV_X1 $T=24940 23400 0 180 $X=24445 $Y=21885
X7075 269 VSS VDD 783 INV_X1 $T=25130 37400 1 0 $X=25015 $Y=35885
X7076 616 VSS VDD 784 INV_X1 $T=25320 15000 0 0 $X=25205 $Y=14885
X7077 953 VSS VDD 280 INV_X1 $T=25510 20600 1 0 $X=25395 $Y=19085
X7078 621 VSS VDD 508 INV_X1 $T=26650 12200 0 0 $X=26535 $Y=12085
X7079 328 VSS VDD 790 INV_X1 $T=27220 26200 1 0 $X=27105 $Y=24685
X7080 954 VSS VDD 310 INV_X1 $T=28550 12200 1 0 $X=28435 $Y=10685
X7081 872 VSS VDD 793 INV_X1 $T=30070 9400 1 0 $X=29955 $Y=7885
X7082 792 VSS VDD 876 INV_X1 $T=30070 26200 1 0 $X=29955 $Y=24685
X7083 631 VSS VDD 900 INV_X1 $T=30830 20600 0 180 $X=30335 $Y=19085
X7084 333 VSS VDD 339 INV_X1 $T=30450 23400 1 0 $X=30335 $Y=21885
X7085 642 VSS VDD 331 INV_X1 $T=30450 29000 1 0 $X=30335 $Y=27485
X7086 873 VSS VDD 938 INV_X1 $T=30640 31800 0 0 $X=30525 $Y=31685
X7087 645 VSS VDD 139 INV_X1 $T=31780 6600 0 180 $X=31285 $Y=5085
X7088 643 VSS VDD 329 INV_X1 $T=31780 37400 1 180 $X=31285 $Y=37285
X7089 646 VSS VDD 341 INV_X1 $T=31780 15000 0 0 $X=31665 $Y=14885
X7090 647 VSS VDD 641 INV_X1 $T=32540 3800 1 180 $X=32045 $Y=3685
X7091 513 VSS VDD 649 INV_X1 $T=32160 40200 0 0 $X=32045 $Y=40085
X7092 800 VSS VDD 656 INV_X1 $T=32350 23400 1 0 $X=32235 $Y=21885
X7093 648 VSS VDD 652 INV_X1 $T=32920 20600 1 0 $X=32805 $Y=19085
X7094 802 VSS VDD 663 INV_X1 $T=33110 9400 1 0 $X=32995 $Y=7885
X7095 653 VSS VDD 356 INV_X1 $T=34060 17800 0 0 $X=33945 $Y=17685
X7096 651 VSS VDD 359 INV_X1 $T=34440 29000 1 0 $X=34325 $Y=27485
X7097 810 VSS VDD 917 INV_X1 $T=35010 15000 0 0 $X=34895 $Y=14885
X7098 669 VSS VDD 665 INV_X1 $T=35580 23400 0 180 $X=35085 $Y=21885
X7099 664 VSS VDD 370 INV_X1 $T=35390 6600 0 0 $X=35275 $Y=6485
X7100 363 VSS VDD 520 INV_X1 $T=35580 34600 0 0 $X=35465 $Y=34485
X7101 378 VSS VDD 364 INV_X1 $T=36150 43000 1 180 $X=35655 $Y=42885
X7102 882 VSS VDD 881 INV_X1 $T=36720 15000 1 180 $X=36225 $Y=14885
X7103 698 VSS VDD 383 INV_X1 $T=36720 37400 1 0 $X=36605 $Y=35885
X7104 883 VSS VDD 404 INV_X1 $T=37860 40200 0 0 $X=37745 $Y=40085
X7105 424 VSS VDD 402 INV_X1 $T=38430 37400 0 180 $X=37935 $Y=35885
X7106 382 VSS VDD 527 INV_X1 $T=38050 43000 1 0 $X=37935 $Y=41485
X7107 885 VSS VDD 436 INV_X1 $T=38240 34600 0 0 $X=38125 $Y=34485
X7108 685 VSS VDD 367 INV_X1 $T=38810 15000 0 180 $X=38315 $Y=13485
X7109 385 VSS VDD 679 INV_X1 $T=38620 23400 0 0 $X=38505 $Y=23285
X7110 409 VSS VDD 912 INV_X1 $T=39190 15000 0 180 $X=38695 $Y=13485
X7111 515 VSS VDD 362 INV_X1 $T=39380 40200 0 180 $X=38885 $Y=38685
X7112 368 VSS VDD 703 INV_X1 $T=39190 26200 0 0 $X=39075 $Y=26085
X7113 318 VSS VDD 428 INV_X1 $T=40140 20600 1 0 $X=40025 $Y=19085
X7114 374 VSS VDD 416 INV_X1 $T=40900 40200 0 180 $X=40405 $Y=38685
X7115 830 VSS VDD 426 INV_X1 $T=41850 29000 0 180 $X=41355 $Y=27485
X7116 371 VSS VDD 419 INV_X1 $T=42230 26200 1 0 $X=42115 $Y=24685
X7117 523 VSS VDD 691 INV_X1 $T=43750 29000 1 180 $X=43255 $Y=28885
X7118 826 VSS VDD 833 INV_X1 $T=44130 40200 0 180 $X=43635 $Y=38685
X7119 707 VSS VDD 448 INV_X1 $T=43940 40200 0 0 $X=43825 $Y=40085
X7120 388 VSS VDD 366 INV_X1 $T=44320 15000 1 0 $X=44205 $Y=13485
X7121 408 VSS VDD 530 INV_X1 $T=44700 20600 1 180 $X=44205 $Y=20485
X7122 710 VSS VDD 468 INV_X1 $T=44320 40200 0 0 $X=44205 $Y=40085
X7123 435 VSS VDD 716 INV_X1 $T=44510 17800 1 0 $X=44395 $Y=16285
X7147 59 VDD 545 541 VSS VSS NOR2_X1 $T=6320 15000 0 0 $X=6205 $Y=14885
X7148 68 VDD 548 52 VSS VSS NOR2_X1 $T=6700 20600 0 0 $X=6585 $Y=20485
X7149 b[29] VDD 546 104 VSS 975 NOR2_X1 $T=7460 1000 1 180 $X=6775 $Y=885
X7150 59 VDD 498 547 VSS VSS NOR2_X1 $T=6890 15000 0 0 $X=6775 $Y=14885
X7151 548 VDD 87 58 VSS VSS NOR2_X1 $T=7270 20600 0 0 $X=7155 $Y=20485
X7152 99 VDD 550 83 VSS VSS NOR2_X1 $T=7460 37400 0 0 $X=7345 $Y=37285
X7153 60 VDD 68 556 VSS VSS NOR2_X1 $T=9360 12200 0 0 $X=9245 $Y=12085
X7154 74 VDD 162 895 VSS VSS NOR2_X1 $T=14490 20600 1 0 $X=14375 $Y=19085
X7155 118 VDD 574 956 VSS VSS NOR2_X1 $T=15250 9400 1 0 $X=15135 $Y=7885
X7156 202 VDD 581 213 VSS VSS NOR2_X1 $T=16580 34600 0 0 $X=16465 $Y=34485
X7157 207 VDD 861 190 VSS VSS NOR2_X1 $T=16960 23400 1 0 $X=16845 $Y=21885
X7158 189 VDD 586 896 VSS VSS NOR2_X1 $T=17530 12200 0 0 $X=17415 $Y=12085
X7159 234 VDD 864 228 VSS VSS NOR2_X1 $T=20190 23400 0 0 $X=20075 $Y=23285
X7160 276 VDD 605 243 VSS VSS NOR2_X1 $T=23990 9400 1 180 $X=23305 $Y=9285
X7161 293 VDD 620 270 VSS VSS NOR2_X1 $T=25510 40200 0 0 $X=25395 $Y=40085
X7162 283 VDD 615 294 VSS VSS NOR2_X1 $T=26650 3800 0 0 $X=26535 $Y=3685
X7163 295 VDD 623 285 VSS VSS NOR2_X1 $T=26650 29000 0 0 $X=26535 $Y=28885
X7164 644 VDD 647 337 VSS 975 NOR2_X1 $T=31590 1000 0 0 $X=31475 $Y=885
X7165 644 VDD 641 645 VSS VSS NOR2_X1 $T=31590 3800 0 0 $X=31475 $Y=3685
X7166 798 VDD 877 357 VSS VSS NOR2_X1 $T=31970 26200 1 0 $X=31855 $Y=24685
X7167 385 VDD 325 522 VSS VSS NOR2_X1 $T=34060 37400 0 180 $X=33375 $Y=35885
X7168 265 VDD 318 809 VSS VSS NOR2_X1 $T=34440 43000 0 0 $X=34325 $Y=42885
X7169 271 VDD 318 662 VSS VSS NOR2_X1 $T=34820 40200 1 0 $X=34705 $Y=38685
X7170 340 VDD 635 369 VSS VSS NOR2_X1 $T=35390 9400 0 0 $X=35275 $Y=9285
X7171 342 VDD 318 811 VSS VSS NOR2_X1 $T=35390 40200 1 0 $X=35275 $Y=38685
X7172 880 VDD 881 812 VSS VSS NOR2_X1 $T=35770 17800 1 0 $X=35655 $Y=16285
X7173 516 VDD 388 424 VSS VSS NOR2_X1 $T=36150 12200 0 0 $X=36035 $Y=12085
X7174 388 VDD 652 471 VSS VSS NOR2_X1 $T=36720 20600 1 180 $X=36035 $Y=20485
X7175 683 VDD 339 344 VSS VSS NOR2_X1 $T=36910 26200 0 180 $X=36225 $Y=24685
X7176 683 VDD 348 346 VSS VSS NOR2_X1 $T=36910 26200 1 0 $X=36795 $Y=24685
X7177 523 VDD 679 351 VSS VSS NOR2_X1 $T=37670 26200 1 180 $X=36985 $Y=26085
X7178 812 VDD 367 397 VSS VSS NOR2_X1 $T=37480 17800 1 0 $X=37365 $Y=16285
X7179 388 VDD 877 472 VSS VSS NOR2_X1 $T=37480 26200 1 0 $X=37365 $Y=24685
X7180 816 VDD 883 886 VSS VSS NOR2_X1 $T=37480 40200 1 0 $X=37365 $Y=38685
X7181 275 VDD 318 910 VSS VSS NOR2_X1 $T=37480 45800 0 0 $X=37365 $Y=45685
X7182 385 VDD 320 674 VSS VSS NOR2_X1 $T=37670 31800 0 0 $X=37555 $Y=31685
X7183 415 VDD 417 403 VSS VSS NOR2_X1 $T=39000 23400 0 0 $X=38885 $Y=23285
X7184 371 VDD 683 377 VSS VSS NOR2_X1 $T=39000 26200 1 0 $X=38885 $Y=24685
X7185 385 VDD 691 514 VSS VSS NOR2_X1 $T=39190 31800 1 0 $X=39075 $Y=30285
X7186 388 VDD 822 470 VSS VSS NOR2_X1 $T=40140 20600 0 180 $X=39455 $Y=19085
X7187 683 VDD 373 412 VSS VSS NOR2_X1 $T=39570 26200 1 0 $X=39455 $Y=24685
X7188 298 VDD 318 958 VSS VSS NOR2_X1 $T=39570 43000 0 0 $X=39455 $Y=42885
X7189 689 VDD 678 824 VSS VSS NOR2_X1 $T=40520 26200 0 0 $X=40405 $Y=26085
X7190 683 VDD 419 694 VSS VSS NOR2_X1 $T=41280 31800 0 0 $X=41165 $Y=31685
X7191 388 VDD 653 478 VSS VSS NOR2_X1 $T=42230 20600 1 0 $X=42115 $Y=19085
X7192 523 VDD 419 831 VSS VSS NOR2_X1 $T=42230 26200 0 0 $X=42115 $Y=26085
X7193 888 VDD 441 887 VSS VSS NOR2_X1 $T=42610 15000 1 0 $X=42495 $Y=13485
X7194 408 VDD 701 834 VSS VSS NOR2_X1 $T=43560 43000 1 180 $X=42875 $Y=42885
X7195 435 VDD 408 432 VSS VSS NOR2_X1 $T=43940 17800 0 180 $X=43255 $Y=16285
X7196 408 VDD 523 466 VSS VSS NOR2_X1 $T=43940 34600 1 0 $X=43825 $Y=33085
X7197 523 VDD 530 705 VSS VSS NOR2_X1 $T=44130 31800 0 0 $X=44015 $Y=31685
X7198 852 44 VSS VDD 36 VSS OR2_X1 $T=4420 40200 0 180 $X=3545 $Y=38685
X7199 536 50 VSS VDD 66 VSS OR2_X1 $T=4610 43000 0 0 $X=4495 $Y=42885
X7200 542 57 VSS VDD 852 VSS OR2_X1 $T=5750 37400 0 180 $X=4875 $Y=35885
X7201 853 b[28] VSS VDD 546 975 OR2_X1 $T=6130 1000 0 0 $X=6015 $Y=885
X7202 858 123 VSS VDD 136 VSS OR2_X1 $T=10500 37400 1 0 $X=10385 $Y=35885
X7203 575 b[27] VSS VDD 853 975 OR2_X1 $T=12020 1000 0 0 $X=11905 $Y=885
X7204 571 146 VSS VDD 858 VSS OR2_X1 $T=12970 34600 1 180 $X=12095 $Y=34485
X7205 743 157 VSS VDD 174 VSS OR2_X1 $T=13920 40200 1 0 $X=13805 $Y=38685
X7206 153 b[26] VSS VDD 575 975 OR2_X1 $T=15440 1000 0 0 $X=15325 $Y=885
X7207 577 176 VSS VDD 861 VSS OR2_X1 $T=16390 29000 1 0 $X=16275 $Y=27485
X7208 584 184 VSS VDD 586 VSS OR2_X1 $T=17340 17800 1 0 $X=17225 $Y=16285
X7209 588 204 VSS VDD 591 VSS OR2_X1 $T=19050 45800 1 0 $X=18935 $Y=44285
X7210 506 212 VSS VDD 594 VSS OR2_X1 $T=20190 17800 0 180 $X=19315 $Y=16285
X7211 760 210 VSS VDD 864 VSS OR2_X1 $T=19430 26200 0 0 $X=19315 $Y=26085
X7212 594 218 VSS VDD 236 VSS OR2_X1 $T=21140 15000 0 180 $X=20265 $Y=13485
X7213 868 256 VSS VDD 610 VSS OR2_X1 $T=24560 31800 1 180 $X=23685 $Y=31685
X7214 601 260 VSS VDD 615 VSS OR2_X1 $T=24750 3800 0 0 $X=24635 $Y=3685
X7215 870 274 VSS VDD 623 VSS OR2_X1 $T=26460 31800 1 180 $X=25585 $Y=31685
X7216 622 271 VSS VDD 625 VSS OR2_X1 $T=25700 40200 1 0 $X=25585 $Y=38685
X7217 640 275 VSS VDD 272 VSS OR2_X1 $T=26460 45800 1 180 $X=25585 $Y=45685
X7218 871 280 VSS VDD 624 VSS OR2_X1 $T=26650 20600 0 0 $X=26535 $Y=20485
X7219 625 290 VSS VDD 321 VSS OR2_X1 $T=27600 43000 1 0 $X=27485 $Y=41485
X7220 628 299 VSS VDD 633 VSS OR2_X1 $T=29120 23400 0 180 $X=28245 $Y=21885
X7221 630 310 VSS VDD 795 VSS OR2_X1 $T=29500 12200 1 0 $X=29385 $Y=10685
X7222 633 314 VSS VDD 311 VSS OR2_X1 $T=29690 20600 1 0 $X=29575 $Y=19085
X7223 638 323 VSS VDD 796 VSS OR2_X1 $T=30640 6600 1 0 $X=30525 $Y=5085
X7224 521 370 VSS VDD 516 VSS OR2_X1 $T=36530 6600 1 180 $X=35655 $Y=6485
X7225 336 385 VSS VDD 681 VSS OR2_X1 $T=36910 31800 0 0 $X=36795 $Y=31685
X7226 324 385 VSS VDD 817 VSS OR2_X1 $T=37480 34600 0 0 $X=37365 $Y=34485
X7227 827 408 VSS VDD 455 VSS OR2_X1 $T=43940 31800 1 0 $X=43825 $Y=30285
X7228 442 408 VSS VDD 944 VSS OR2_X1 $T=44130 23400 0 0 $X=44015 $Y=23285
X7238 9 8 a[29] 850 VDD VSS 17 975 FA_X1 $T=1000 1000 0 0 $X=885 $Y=885
X7239 537 9 a[30] 851 VDD VSS 849 VSS FA_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X7240 8 48 a[28] 538 VDD VSS 543 VSS FA_X1 $T=4040 3800 0 0 $X=3925 $Y=3685
X7241 48 88 a[27] 857 VDD VSS 97 VSS FA_X1 $T=7080 3800 0 0 $X=6965 $Y=3685
X7242 124 114 a[25] 855 VDD VSS 497 VSS FA_X1 $T=10690 6600 0 180 $X=7535 $Y=5085
X7243 88 124 a[26] 860 VDD VSS 105 VSS FA_X1 $T=10120 3800 0 0 $X=10005 $Y=3685
X7244 114 130 a[24] 750 VDD VSS 109 VSS FA_X1 $T=10500 6600 0 0 $X=10385 $Y=6485
X7245 803 350 932 379 VDD VSS 360 VSS FA_X1 $T=33300 3800 0 0 $X=33185 $Y=3685
X7246 350 921 413 379 VDD VSS 410 VSS FA_X1 $T=41850 6600 0 180 $X=38695 $Y=5085
X7247 430 406 465 887 VDD VSS 457 VSS FA_X1 $T=38810 6600 0 0 $X=38695 $Y=6485
X7248 921 430 709 890 VDD VSS 454 VSS FA_X1 $T=41850 3800 0 0 $X=41735 $Y=3685
X7249 406 450 463 891 VDD VSS 477 VSS FA_X1 $T=43750 9400 1 0 $X=43635 $Y=7885
X7250 450 451 439 892 VDD VSS 485 VSS FA_X1 $T=43750 12200 0 0 $X=43635 $Y=12085
X7265 117 17 35 539 VSS VDD AOI21_X1 $T=2900 9400 0 180 $X=2025 $Y=7885
X7266 117 97 64 553 VSS VDD AOI21_X1 $T=7840 9400 1 0 $X=7725 $Y=7885
X7267 560 155 169 895 VSS VDD AOI21_X1 $T=13730 20600 1 0 $X=13615 $Y=19085
X7268 894 175 276 755 VSS VDD AOI21_X1 $T=15820 9400 0 0 $X=15705 $Y=9285
X7269 915 179 273 755 VSS VDD AOI21_X1 $T=17340 9400 1 180 $X=16465 $Y=9285
X7270 900 333 822 957 VSS VDD AOI21_X1 $T=29690 17800 0 0 $X=29575 $Y=17685
X7271 903 329 901 634 VSS VDD AOI21_X1 $T=30640 37400 0 0 $X=30525 $Y=37285
X7272 874 331 798 511 VSS VDD AOI21_X1 $T=30830 29000 1 0 $X=30715 $Y=27485
X7273 876 333 877 639 VSS VDD AOI21_X1 $T=31210 26200 1 0 $X=31095 $Y=24685
X7274 341 333 653 797 VSS VDD AOI21_X1 $T=32920 17800 1 0 $X=32805 $Y=16285
X7275 342 339 372 939 VSS VDD AOI21_X1 $T=34820 40200 0 180 $X=33945 $Y=38685
X7276 822 356 880 917 VSS VDD AOI21_X1 $T=34250 17800 1 0 $X=34135 $Y=16285
X7277 297 339 391 916 VSS VDD AOI21_X1 $T=35390 45800 0 180 $X=34515 $Y=44285
X7278 318 362 343 809 VSS VDD AOI21_X1 $T=35580 40200 1 180 $X=34705 $Y=40085
X7279 819 364 878 375 VSS VDD AOI21_X1 $T=35010 43000 0 0 $X=34895 $Y=42885
X7280 371 368 908 814 VSS VDD AOI21_X1 $T=36340 26200 1 180 $X=35465 $Y=26085
X7281 318 372 820 662 VSS VDD AOI21_X1 $T=36720 40200 0 180 $X=35845 $Y=38685
X7282 657 377 437 908 VSS VDD AOI21_X1 $T=36150 23400 1 0 $X=36035 $Y=21885
X7283 371 380 909 918 VSS VDD AOI21_X1 $T=36340 26200 0 0 $X=36225 $Y=26085
X7284 385 383 885 522 VSS VDD AOI21_X1 $T=37480 34600 1 180 $X=36605 $Y=34485
X7285 318 383 883 811 VSS VDD AOI21_X1 $T=37480 40200 0 180 $X=36605 $Y=38685
X7286 377 389 920 909 VSS VDD AOI21_X1 $T=36910 23400 1 0 $X=36795 $Y=21885
X7287 318 391 375 910 VSS VDD AOI21_X1 $T=38050 45800 0 180 $X=37175 $Y=44285
X7288 393 395 948 398 VSS VDD AOI21_X1 $T=37670 23400 1 0 $X=37555 $Y=21885
X7289 816 404 884 820 VSS VDD AOI21_X1 $T=39760 40200 1 180 $X=38885 $Y=40085
X7290 429 412 386 424 VSS VDD AOI21_X1 $T=39570 37400 1 0 $X=39455 $Y=35885
X7291 318 416 382 958 VSS VDD AOI21_X1 $T=40900 43000 1 180 $X=40025 $Y=42885
X7292 385 416 696 674 VSS VDD AOI21_X1 $T=40520 31800 0 0 $X=40405 $Y=31685
X7293 419 414 431 824 VSS VDD AOI21_X1 $T=40710 23400 1 0 $X=40595 $Y=21885
X7294 387 433 889 834 VSS VDD AOI21_X1 $T=42230 43000 0 0 $X=42115 $Y=42885
X7295 419 432 888 679 VSS VDD AOI21_X1 $T=44130 17800 1 180 $X=43255 $Y=17685
X7333 536 51 VSS VDD 100 AND2_X1 $T=4610 45800 0 0 $X=4495 $Y=45685
X7334 498 59 VSS VDD 122 AND2_X1 $T=5560 15000 0 0 $X=5445 $Y=14885
X7335 542 63 VSS VDD 75 AND2_X1 $T=5750 34600 0 0 $X=5635 $Y=34485
X7336 550 91 VSS VDD 92 AND2_X1 $T=7460 40200 0 0 $X=7345 $Y=40085
X7337 574 117 VSS VDD 502 AND2_X1 $T=10120 9400 1 0 $X=10005 $Y=7885
X7338 743 141 VSS VDD 144 AND2_X1 $T=11830 40200 1 0 $X=11715 $Y=38685
X7339 924 142 VSS VDD 561 AND2_X1 $T=11830 43000 0 0 $X=11715 $Y=42885
X7340 74 111 VSS VDD 565 AND2_X1 $T=12210 12200 0 0 $X=12095 $Y=12085
X7341 153 151 VSS VDD 855 AND2_X1 $T=13920 3800 1 180 $X=13045 $Y=3685
X7342 571 160 VSS VDD 165 AND2_X1 $T=14490 34600 0 0 $X=14375 $Y=34485
X7343 581 177 VSS VDD 183 AND2_X1 $T=16390 40200 1 0 $X=16275 $Y=38685
X7344 589 203 VSS VDD 588 AND2_X1 $T=19430 45800 1 180 $X=18555 $Y=45685
X7345 772 216 VSS VDD 768 AND2_X1 $T=20760 43000 0 180 $X=19885 $Y=41485
X7346 768 231 VSS VDD 600 AND2_X1 $T=21140 45800 1 0 $X=21025 $Y=44285
X7347 600 233 VSS VDD 589 AND2_X1 $T=21900 45800 1 180 $X=21025 $Y=45685
X7348 602 244 VSS VDD 780 AND2_X1 $T=23040 29000 1 180 $X=22165 $Y=28885
X7349 605 245 VSS VDD 249 AND2_X1 $T=22660 12200 1 0 $X=22545 $Y=10685
X7350 591 251 VSS VDD 607 AND2_X1 $T=23990 45800 0 180 $X=23115 $Y=44285
X7351 607 253 VSS VDD 611 AND2_X1 $T=23610 43000 0 0 $X=23495 $Y=42885
X7352 613 261 VSS VDD 614 AND2_X1 $T=24750 17800 0 0 $X=24635 $Y=17685
X7353 507 262 VSS VDD 785 AND2_X1 $T=24940 29000 1 0 $X=24825 $Y=27485
X7354 786 277 VSS VDD 871 AND2_X1 $T=26270 23400 1 0 $X=26155 $Y=21885
X7355 620 278 VSS VDD 306 AND2_X1 $T=26270 43000 0 0 $X=26155 $Y=42885
X7356 622 281 VSS VDD 338 AND2_X1 $T=26650 37400 0 0 $X=26535 $Y=37285
X7357 624 284 VSS VDD 787 AND2_X1 $T=27600 20600 0 180 $X=26725 $Y=19085
X7358 787 286 VSS VDD 791 AND2_X1 $T=27220 17800 1 0 $X=27105 $Y=16285
X7359 791 291 VSS VDD 629 AND2_X1 $T=27790 15000 1 0 $X=27675 $Y=13485
X7360 635 952 VSS VDD 646 AND2_X1 $T=30070 15000 0 0 $X=29955 $Y=14885
X7361 640 326 VSS VDD 384 AND2_X1 $T=30640 45800 0 0 $X=30525 $Y=45685
X7362 795 330 VSS VDD 655 AND2_X1 $T=31020 12200 1 0 $X=30905 $Y=10685
X7363 338 348 VSS VDD 939 AND2_X1 $T=33300 40200 1 0 $X=33185 $Y=38685
X7364 655 349 VSS VDD 806 AND2_X1 $T=33490 9400 0 0 $X=33375 $Y=9285
X7365 384 348 VSS VDD 916 AND2_X1 $T=34060 45800 0 0 $X=33945 $Y=45685
X7366 806 365 VSS VDD 668 AND2_X1 $T=35390 9400 1 0 $X=35275 $Y=7885
X7367 668 392 VSS VDD 521 AND2_X1 $T=38050 9400 0 180 $X=37175 $Y=7885
X7368 816 438 VSS VDD sum[0] AND2_X1 $T=42800 29000 1 0 $X=42685 $Y=27485
X7380 541 VSS 60 68 VDD 128 NAND3_X1 $T=7840 17800 1 0 $X=7725 $Y=16285
X7381 118 VSS 574 108 VDD 915 NAND3_X1 $T=15820 12200 1 0 $X=15705 $Y=10685
X7382 371 VSS 381 679 VDD 699 NAND3_X1 $T=43180 34600 1 180 $X=42305 $Y=34485
X7481 85 49 VDD 58 60 61 VSS 87 112 AOI222_X1 $T=4990 20600 1 0 $X=4875 $Y=19085
X7482 58 115 VDD 81 85 87 VSS 72 107 AOI222_X1 $T=6510 26200 1 0 $X=6395 $Y=24685
X7483 58 79 VDD 102 85 87 VSS 730 126 AOI222_X1 $T=8030 26200 1 0 $X=7915 $Y=24685
X7484 58 129 VDD 106 85 87 VSS 98 134 AOI222_X1 $T=8410 20600 1 0 $X=8295 $Y=19085
X7485 52 140 VDD 85 115 111 VSS 119 156 AOI222_X1 $T=10880 23400 0 180 $X=9245 $Y=21885
X7486 81 111 VDD 85 119 122 VSS 563 147 AOI222_X1 $T=9550 23400 0 0 $X=9435 $Y=23285
X7487 106 111 VDD 85 125 122 VSS 133 154 AOI222_X1 $T=9930 20600 1 0 $X=9815 $Y=19085
X7488 52 110 VDD 85 79 111 VSS 727 163 AOI222_X1 $T=10880 23400 1 0 $X=10765 $Y=21885
X7489 52 118 VDD 85 129 111 VSS 125 162 AOI222_X1 $T=11450 17800 0 0 $X=11335 $Y=17685
X7490 727 85 VDD 111 102 122 VSS 155 145 AOI222_X1 $T=12780 26200 1 0 $X=12665 $Y=24685
X7491 792 344 VDD 346 328 351 VSS 515 380 AOI222_X1 $T=32920 26200 0 0 $X=32805 $Y=26085
X7492 409 428 VDD 420 421 424 VSS 394 828 AOI222_X1 $T=40330 15000 0 0 $X=40215 $Y=14885
X7493 394 428 VDD 429 421 424 VSS 355 721 AOI222_X1 $T=41280 17800 0 0 $X=41165 $Y=17685
X7494 728 VDD 534 893 VSS 741 NOR3_X1 $T=5560 9400 0 180 $X=4685 $Y=7885
X7495 68 VDD 59 498 VSS 551 NOR3_X1 $T=4990 15000 1 0 $X=4875 $Y=13485
X7496 74 VDD 59 545 VSS 567 NOR3_X1 $T=9930 15000 1 0 $X=9815 $Y=13485
X7497 545 VDD 59 108 VSS 560 NOR3_X1 $T=10120 15000 0 0 $X=10005 $Y=14885
X7498 74 VDD 574 755 VSS 208 NOR3_X1 $T=15820 9400 1 0 $X=15705 $Y=7885
X7499 214 VDD 207 861 VSS 186 NOR3_X1 $T=16960 23400 0 180 $X=16085 $Y=21885
X7500 74 VDD 956 755 VSS 225 NOR3_X1 $T=16580 9400 1 0 $X=16465 $Y=7885
X7501 196 VDD 189 586 VSS 223 NOR3_X1 $T=18860 12200 1 180 $X=17985 $Y=12085
X7502 273 VDD 276 605 VSS 226 NOR3_X1 $T=20000 9400 0 0 $X=19885 $Y=9285
X7503 164 VDD 234 864 VSS 863 NOR3_X1 $T=20760 20600 1 180 $X=19885 $Y=20485
X7504 305 VDD 295 623 VSS 304 NOR3_X1 $T=27030 29000 1 0 $X=26915 $Y=27485
X7505 317 VDD 283 615 VSS 323 NOR3_X1 $T=27980 3800 1 180 $X=27105 $Y=3685
X7506 875 VDD 873 642 VSS 512 NOR3_X1 $T=30830 31800 1 0 $X=30715 $Y=30285
X7507 902 VDD 634 332 VSS 875 NOR3_X1 $T=30830 34600 0 0 $X=30715 $Y=34485
X7508 940 VDD 513 643 VSS 902 NOR3_X1 $T=32160 40200 1 180 $X=31285 $Y=40085
X7509 512 VDD 511 877 VSS 801 NOR3_X1 $T=32160 26200 0 0 $X=32045 $Y=26085
X7510 801 VDD 656 652 VSS 904 NOR3_X1 $T=32730 20600 0 0 $X=32615 $Y=20485
X7511 904 VDD 822 653 VSS 805 NOR3_X1 $T=33300 17800 0 0 $X=33185 $Y=17685
X7512 805 VDD 917 881 VSS 818 NOR3_X1 $T=35010 17800 1 0 $X=34895 $Y=16285
X7513 813 VDD 375 343 VSS 940 NOR3_X1 $T=36150 43000 0 180 $X=35275 $Y=41485
X7514 680 VDD 382 378 VSS 813 NOR3_X1 $T=38050 43000 0 180 $X=37175 $Y=41485
X7515 886 VDD 820 399 VSS 680 NOR3_X1 $T=38240 40200 0 0 $X=38125 $Y=40085
X7516 355 VDD 340 635 VSS 411 NOR3_X1 $T=38620 12200 1 0 $X=38505 $Y=10685
X7517 714 VDD 683 373 VSS 667 NOR3_X1 $T=39570 29000 0 0 $X=39455 $Y=28885
X7518 385 VDD 435 373 VSS 441 NOR3_X1 $T=40520 17800 0 0 $X=40405 $Y=17685
X7519 530 VDD 371 683 VSS 433 NOR3_X1 $T=41090 34600 0 0 $X=40975 $Y=34485
X7520 558 500 VSS 123 172 127 VDD OAI22_X1 $T=9930 31800 0 0 $X=9815 $Y=31685
X7521 558 127 VSS 132 172 749 VDD OAI22_X1 $T=10880 31800 0 0 $X=10765 $Y=31685
X7522 558 742 VSS 173 172 745 VDD OAI22_X1 $T=11070 31800 1 0 $X=10955 $Y=30285
X7523 558 745 VSS 146 172 500 VDD OAI22_X1 $T=11830 31800 0 0 $X=11715 $Y=31685
X7524 558 749 VSS 135 172 928 VDD OAI22_X1 $T=12780 31800 0 0 $X=12665 $Y=31685
X7525 558 740 VSS 148 172 927 VDD OAI22_X1 $T=13160 29000 0 0 $X=13045 $Y=28885
X7526 172 742 VSS 150 558 927 VDD OAI22_X1 $T=13350 31800 1 0 $X=13235 $Y=30285
X7527 558 928 VSS 157 172 570 VDD OAI22_X1 $T=13730 31800 0 0 $X=13615 $Y=31685
X7528 172 752 VSS 166 570 558 VDD OAI22_X1 $T=14300 31800 1 0 $X=14185 $Y=30285
X7529 566 172 VSS 246 572 558 VDD OAI22_X1 $T=16010 17800 1 180 $X=14945 $Y=17685
X7530 172 572 VSS 164 169 558 VDD OAI22_X1 $T=15060 20600 1 0 $X=14945 $Y=19085
X7531 558 566 VSS 212 172 753 VDD OAI22_X1 $T=16200 17800 0 180 $X=15135 $Y=16285
X7532 752 558 VSS 170 754 172 VDD OAI22_X1 $T=15250 31800 1 0 $X=15135 $Y=30285
X7533 558 753 VSS 218 172 576 VDD OAI22_X1 $T=15440 15000 0 0 $X=15325 $Y=14885
X7534 558 576 VSS 232 929 172 VDD OAI22_X1 $T=15630 15000 1 0 $X=15515 $Y=13485
X7535 172 580 VSS 210 930 558 VDD OAI22_X1 $T=16580 26200 0 180 $X=15515 $Y=24685
X7536 558 751 VSS 230 172 930 VDD OAI22_X1 $T=15820 26200 0 0 $X=15705 $Y=26085
X7537 172 751 VSS 202 754 558 VDD OAI22_X1 $T=17150 31800 0 180 $X=16085 $Y=30285
X7538 578 172 VSS 227 929 558 VDD OAI22_X1 $T=16580 12200 0 0 $X=16465 $Y=12085
X7539 580 558 VSS 234 169 172 VDD OAI22_X1 $T=16580 20600 0 0 $X=16465 $Y=20485
X7540 299 318 VSS 639 328 335 VDD OAI22_X1 $T=30260 23400 0 0 $X=30145 $Y=23285
X7541 313 318 VSS 957 312 335 VDD OAI22_X1 $T=30450 17800 0 0 $X=30335 $Y=17685
X7542 340 318 VSS 797 313 335 VDD OAI22_X1 $T=32350 15000 0 180 $X=31285 $Y=13485
X7543 274 318 VSS 474 402 324 VDD OAI22_X1 $T=31590 34600 0 0 $X=31475 $Y=34485
X7544 295 318 VSS 483 402 320 VDD OAI22_X1 $T=31780 31800 0 0 $X=31665 $Y=31685
X7545 267 318 VSS 476 402 336 VDD OAI22_X1 $T=32350 45800 1 0 $X=32235 $Y=44285
X7546 269 318 VSS 484 402 308 VDD OAI22_X1 $T=32540 37400 1 0 $X=32425 $Y=35885
X7547 293 318 VSS 475 402 325 VDD OAI22_X1 $T=32540 40200 0 0 $X=32425 $Y=40085
X7548 328 318 VSS 482 402 334 VDD OAI22_X1 $T=33490 29000 1 0 $X=33375 $Y=27485
X7549 305 318 VSS 473 402 322 VDD OAI22_X1 $T=33490 29000 0 0 $X=33375 $Y=28885
X7550 265 318 VSS 456 402 515 VDD OAI22_X1 $T=38050 45800 0 0 $X=37935 $Y=45685
X7551 362 684 VSS 682 371 688 VDD OAI22_X1 $T=40140 34600 1 180 $X=39075 $Y=34485
X7552 688 689 VSS 462 371 380 VDD OAI22_X1 $T=40520 26200 1 180 $X=39455 $Y=26085
X7553 391 684 VSS 460 692 371 VDD OAI22_X1 $T=40140 34600 0 0 $X=40025 $Y=34485
X7554 297 318 VSS 434 402 381 VDD OAI22_X1 $T=40140 45800 0 0 $X=40025 $Y=45685
X7555 689 692 VSS 445 678 832 VDD OAI22_X1 $T=40900 29000 0 0 $X=40785 $Y=28885
X7556 416 684 VSS 825 427 371 VDD OAI22_X1 $T=40900 34600 1 0 $X=40785 $Y=33085
X7557 275 318 VSS 444 402 815 VDD OAI22_X1 $T=40900 45800 1 0 $X=40785 $Y=44285
X7599 636 339 VSS 318 314 335 VDD 299 800 OAI222_X1 $T=30830 23400 1 0 $X=30715 $Y=21885
X7600 632 339 VSS 318 312 335 VDD 314 648 OAI222_X1 $T=31210 20600 0 0 $X=31095 $Y=20485
X7601 345 339 VSS 318 355 335 VDD 340 810 OAI222_X1 $T=33680 15000 1 0 $X=33565 $Y=13485
X7602 376 339 VSS 318 394 335 VDD 355 882 OAI222_X1 $T=38810 15000 1 180 $X=37175 $Y=14885
X7603 390 339 VSS 318 409 335 VDD 394 685 OAI222_X1 $T=38810 15000 0 0 $X=38695 $Y=14885
X7604 225 VDD 273 276 605 195 VSS NOR4_X1 $T=18670 9400 1 0 $X=18555 $Y=7885
X7605 873 VDD 642 511 877 659 VSS NOR4_X1 $T=31210 29000 0 0 $X=31095 $Y=28885
X7606 513 VDD 643 634 332 347 VSS NOR4_X1 $T=32540 37400 0 180 $X=31475 $Y=35885
X7607 656 VDD 652 822 653 361 VSS NOR4_X1 $T=33490 20600 0 0 $X=33375 $Y=20485
X7608 652 VDD 653 881 400 661 VSS NOR4_X1 $T=35010 20600 1 0 $X=34895 $Y=19085
X7609 917 VDD 881 367 400 669 VSS NOR4_X1 $T=35390 17800 0 0 $X=35275 $Y=17685
X7610 394 VDD 355 340 635 407 VSS NOR4_X1 $T=37860 9400 0 0 $X=37745 $Y=9285
X7611 816 VDD 883 820 399 524 VSS NOR4_X1 $T=38050 40200 1 0 $X=37935 $Y=38685
X7612 545 111 59 68 VSS VDD NOR3_X2 $T=4230 12200 1 0 $X=4115 $Y=10685
X7613 87 85 59 545 VSS VDD NOR3_X2 $T=7840 15000 0 0 $X=7725 $Y=14885
X7614 400 408 367 818 VSS VDD NOR3_X2 $T=39380 17800 0 180 $X=37935 $Y=16285
X7615 VDD 42 70 36 VSS VSS XOR2_X1 $T=2140 45800 1 180 $X=885 $Y=45685
X7616 VDD 17 534 539 VSS VSS XOR2_X1 $T=2330 6600 0 0 $X=2215 $Y=6485
X7617 VDD b[29] 850 546 VSS 975 XOR2_X1 $T=5180 1000 1 180 $X=3925 $Y=885
X7618 VDD 44 73 852 VSS VSS XOR2_X1 $T=4420 40200 1 0 $X=4305 $Y=38685
X7619 VDD b[28] 538 853 VSS VSS XOR2_X1 $T=6320 3800 0 180 $X=5065 $Y=2285
X7620 VDD 99 90 550 VSS VSS XOR2_X1 $T=6320 37400 0 0 $X=6205 $Y=37285
X7621 VDD 105 59 732 VSS VSS XOR2_X1 $T=7270 12200 1 0 $X=7155 $Y=10685
X7622 VDD 56 131 53 VSS VSS XOR2_X1 $T=8220 34600 1 0 $X=8105 $Y=33085
X7623 VDD 132 138 136 VSS VSS XOR2_X1 $T=8790 40200 1 0 $X=8675 $Y=38685
X7624 VDD b[27] 857 575 VSS 975 XOR2_X1 $T=12020 1000 1 180 $X=10765 $Y=885
X7625 VDD 142 216 924 VSS VSS XOR2_X1 $T=11450 43000 1 0 $X=11335 $Y=41485
X7626 VDD 561 231 738 VSS VSS XOR2_X1 $T=12590 43000 0 0 $X=12475 $Y=42885
X7627 VDD 564 233 562 VSS VSS XOR2_X1 $T=12970 45800 0 0 $X=12855 $Y=45685
X7628 VDD b[24] 750 b[23] VSS VSS XOR2_X1 $T=14490 6600 0 180 $X=13235 $Y=5085
X7629 VDD 157 171 743 VSS VSS XOR2_X1 $T=13350 40200 0 0 $X=13235 $Y=40085
X7630 VDD b[26] 860 153 VSS VSS XOR2_X1 $T=15630 3800 0 180 $X=14375 $Y=2285
X7631 VDD 166 167 174 VSS VSS XOR2_X1 $T=14490 40200 0 0 $X=14375 $Y=40085
X7632 VDD 756 573 926 VSS VSS XOR2_X1 $T=14490 45800 1 0 $X=14375 $Y=44285
X7633 VDD 202 194 581 VSS VSS XOR2_X1 $T=16010 37400 1 0 $X=15895 $Y=35885
X7634 VDD 184 209 584 VSS VSS XOR2_X1 $T=17340 17800 0 180 $X=16085 $Y=16285
X7635 VDD 582 203 573 VSS VSS XOR2_X1 $T=17530 45800 0 0 $X=17415 $Y=45685
X7636 VDD 189 197 586 VSS VSS XOR2_X1 $T=18100 15000 1 0 $X=17985 $Y=13485
X7637 VDD 232 240 236 VSS VSS XOR2_X1 $T=19240 15000 1 0 $X=19125 $Y=13485
X7638 VDD 589 275 203 VSS VSS XOR2_X1 $T=19430 45800 0 0 $X=19315 $Y=45685
X7639 VDD 766 255 759 VSS VSS XOR2_X1 $T=20190 34600 1 0 $X=20075 $Y=33085
X7640 VDD 212 241 506 VSS VSS XOR2_X1 $T=20760 17800 0 0 $X=20645 $Y=17685
X7641 VDD 774 599 898 VSS VSS XOR2_X1 $T=20760 31800 0 0 $X=20645 $Y=31685
X7642 VDD 772 290 216 VSS VSS XOR2_X1 $T=20760 43000 1 0 $X=20645 $Y=41485
X7643 VDD 768 298 231 VSS VSS XOR2_X1 $T=20760 43000 0 0 $X=20645 $Y=42885
X7644 VDD 276 266 605 VSS VSS XOR2_X1 $T=22280 9400 0 0 $X=22165 $Y=9285
X7645 VDD 780 262 777 VSS VSS XOR2_X1 $T=22280 29000 1 0 $X=22165 $Y=27485
X7646 VDD 771 342 762 VSS VSS XOR2_X1 $T=22280 37400 1 0 $X=22165 $Y=35885
X7647 VDD 595 271 592 VSS VSS XOR2_X1 $T=22280 37400 0 0 $X=22165 $Y=37285
X7648 VDD 600 297 233 VSS VSS XOR2_X1 $T=22280 45800 0 0 $X=22165 $Y=45685
X7649 VDD 775 934 608 VSS VSS XOR2_X1 $T=23420 20600 1 0 $X=23305 $Y=19085
X7650 VDD 778 269 254 VSS VSS XOR2_X1 $T=23420 37400 1 0 $X=23305 $Y=35885
X7651 VDD 591 265 251 VSS VSS XOR2_X1 $T=23420 45800 0 0 $X=23305 $Y=45685
X7652 VDD 261 284 613 VSS VSS XOR2_X1 $T=23610 17800 0 0 $X=23495 $Y=17685
X7653 VDD 610 274 259 VSS VSS XOR2_X1 $T=23800 31800 1 0 $X=23685 $Y=30285
X7654 VDD 782 277 934 VSS VSS XOR2_X1 $T=24180 20600 0 0 $X=24065 $Y=20485
X7655 VDD 265 301 272 VSS VSS XOR2_X1 $T=24560 45800 0 0 $X=24445 $Y=45685
X7656 VDD 271 319 622 VSS VSS XOR2_X1 $T=24750 37400 0 0 $X=24635 $Y=37285
X7657 VDD 614 286 936 VSS VSS XOR2_X1 $T=24940 17800 1 0 $X=24825 $Y=16285
X7658 VDD 507 295 262 VSS VSS XOR2_X1 $T=24940 29000 0 0 $X=24825 $Y=28885
X7659 VDD 283 279 615 VSS VSS XOR2_X1 $T=25510 3800 0 0 $X=25395 $Y=3685
X7660 VDD 786 328 277 VSS VSS XOR2_X1 $T=25510 23400 0 0 $X=25395 $Y=23285
X7661 VDD 255 302 257 VSS VSS XOR2_X1 $T=25510 34600 1 0 $X=25395 $Y=33085
X7662 VDD 784 291 781 VSS VSS XOR2_X1 $T=25700 15000 1 0 $X=25585 $Y=13485
X7663 VDD 785 305 268 VSS VSS XOR2_X1 $T=25700 26200 0 0 $X=25585 $Y=26085
X7664 VDD 293 288 620 VSS VSS XOR2_X1 $T=26460 43000 1 0 $X=26345 $Y=41485
X7665 VDD 787 314 286 VSS VSS XOR2_X1 $T=27030 17800 0 0 $X=26915 $Y=17685
X7666 VDD 295 300 623 VSS VSS XOR2_X1 $T=27030 31800 1 0 $X=26915 $Y=30285
X7667 VDD 791 312 291 VSS VSS XOR2_X1 $T=27220 15000 0 0 $X=27105 $Y=14885
X7668 VDD 624 299 284 VSS VSS XOR2_X1 $T=27410 20600 0 0 $X=27295 $Y=20485
X7669 VDD 290 316 625 VSS VSS XOR2_X1 $T=27980 40200 1 0 $X=27865 $Y=38685
X7670 VDD 629 313 303 VSS VSS XOR2_X1 $T=28550 15000 1 0 $X=28435 $Y=13485
X7671 VDD 312 631 311 VSS VSS XOR2_X1 $T=28550 20600 1 0 $X=28435 $Y=19085
X7672 VDD 314 632 633 VSS VSS XOR2_X1 $T=28550 20600 0 0 $X=28435 $Y=20485
X7673 VDD 299 636 628 VSS VSS XOR2_X1 $T=29120 23400 0 0 $X=29005 $Y=23285
X7674 VDD 275 794 640 VSS VSS XOR2_X1 $T=29500 45800 0 0 $X=29385 $Y=45685
X7675 VDD 598 509 637 VSS VSS XOR2_X1 $T=29690 6600 0 0 $X=29575 $Y=6485
X7676 VDD 298 352 321 VSS VSS XOR2_X1 $T=29880 43000 0 0 $X=29765 $Y=42885
X7677 VDD 627 349 789 VSS VSS XOR2_X1 $T=30070 9400 0 0 $X=29955 $Y=9285
X7678 VDD 795 340 330 VSS VSS XOR2_X1 $T=31210 9400 0 0 $X=31095 $Y=9285
X7679 VDD 793 365 509 VSS VSS XOR2_X1 $T=31970 9400 1 0 $X=31855 $Y=7885
X7680 VDD 340 345 635 VSS VSS XOR2_X1 $T=31970 12200 0 0 $X=31855 $Y=12085
X7681 VDD 655 355 349 VSS VSS XOR2_X1 $T=33490 9400 1 180 $X=32235 $Y=9285
X7682 VDD 663 392 804 VSS VSS XOR2_X1 $T=34250 9400 1 0 $X=34135 $Y=7885
X7683 VDD 806 394 365 VSS VSS XOR2_X1 $T=34250 9400 0 0 $X=34135 $Y=9285
X7684 VDD 668 409 392 VSS VSS XOR2_X1 $T=38050 9400 1 0 $X=37935 $Y=7885
X7730 492 VSS VDD 117 CLKBUF_X1 $T=2330 9400 0 0 $X=2215 $Y=9285
X7731 492 VSS VDD 37 CLKBUF_X1 $T=3470 9400 0 0 $X=3355 $Y=9285
X7732 333 VSS VDD 348 CLKBUF_X1 $T=35200 15000 1 0 $X=35085 $Y=13485
X7733 518 VDD 659 385 347 VSS AOI21_X2 $T=32920 31800 1 0 $X=32805 $Y=30285
X7734 665 VDD 358 371 361 VSS AOI21_X2 $T=35770 23400 1 180 $X=34325 $Y=23285
X7735 VSS VDD 123 116 858 ICV_33 $T=8220 37400 1 0 $X=8105 $Y=35885
X7736 VSS VDD 176 187 577 ICV_33 $T=14110 29000 0 0 $X=13995 $Y=28885
X7737 VSS VDD 150 181 148 ICV_33 $T=14680 31800 0 0 $X=14565 $Y=31685
X7738 VSS VDD 758 253 587 ICV_33 $T=18480 43000 0 0 $X=18365 $Y=42885
X7739 VSS VDD 260 263 601 ICV_33 $T=22280 6600 0 0 $X=22165 $Y=6485
X7740 VSS VDD 611 293 250 ICV_33 $T=22280 40200 0 0 $X=22165 $Y=40085
X7741 VSS VDD 607 267 253 ICV_33 $T=22280 43000 1 0 $X=22165 $Y=41485
X7742 VSS VDD 808 804 796 ICV_33 $T=31780 6600 1 0 $X=31665 $Y=5085
X7751 36 42 45 VSS VDD 536 VSS OR3_X1 $T=3660 43000 0 0 $X=3545 $Y=42885
X7752 86 56 53 VSS VDD 542 VSS OR3_X1 $T=5750 34600 0 180 $X=4685 $Y=33085
X7753 66 76 80 VSS VDD 550 VSS OR3_X1 $T=6510 43000 1 0 $X=6395 $Y=41485
X7754 136 132 135 VSS VDD 743 VSS OR3_X1 $T=11070 37400 0 0 $X=10955 $Y=37285
X7755 173 150 148 VSS VDD 571 VSS OR3_X1 $T=13730 34600 0 180 $X=12665 $Y=33085
X7756 b[25] b[24] b[23] VSS VDD 153 975 OR3_X1 $T=14490 1000 0 0 $X=14375 $Y=885
X7757 174 166 170 VSS VDD 581 VSS OR3_X1 $T=15250 37400 0 0 $X=15135 $Y=37285
X7758 236 232 227 VSS VDD 605 VSS OR3_X1 $T=21900 12200 0 180 $X=20835 $Y=10685
X7759 342 255 257 VSS VDD 622 VSS OR3_X1 $T=23800 37400 0 0 $X=23685 $Y=37285
X7760 272 265 267 VSS VDD 620 VSS OR3_X1 $T=25320 43000 0 0 $X=25205 $Y=42885
X7761 321 298 297 VSS VDD 640 VSS OR3_X1 $T=28930 45800 0 180 $X=27865 $Y=44285
X7762 311 312 313 VSS VDD 635 VSS OR3_X1 $T=29500 17800 1 0 $X=29385 $Y=16285
X7763 a[2] 37 b[2] VSS VDD 86 b[2] 18 a[2] 725 VSS ICV_35 $T=1000 12200 0 0 $X=885 $Y=12085
X7764 b[5] 18 a[5] VSS VDD 726 b[17] 18 a[17] 115 VSS ICV_35 $T=2330 23400 1 0 $X=2215 $Y=21885
X7765 a[12] 37 b[12] VSS VDD 176 b[12] 18 a[12] 727 VSS ICV_35 $T=2330 26200 0 0 $X=2215 $Y=26085
X7766 b[13] 18 a[13] VSS VDD 119 a[13] 37 b[13] 207 VSS ICV_35 $T=3660 23400 0 0 $X=3545 $Y=23285
X7767 b[18] 18 a[18] VSS VDD 129 a[18] 37 b[18] 196 VSS ICV_35 $T=18100 3800 0 0 $X=17985 $Y=3685
X7768 a[19] 37 b[19] VSS VDD 247 b[22] 18 a[22] 118 VSS ICV_35 $T=19240 3800 1 0 $X=19125 $Y=2285
X7769 206 638 214 VSS VDD 609 219 139 164 933 VSS ICV_35 $T=19240 23400 1 0 $X=19125 $Y=21885
X7770 b[21] 18 a[21] VSS VDD 140 a[21] 37 b[21] 283 975 ICV_35 $T=23040 1000 0 0 $X=22925 $Y=885
X7771 295 333 300 VSS VDD 322 295 318 320 873 VSS ICV_35 $T=28170 31800 1 0 $X=28055 $Y=30285
X7772 b[31] 18 a[31] VSS VDD 647 a[31] 37 b[31] 644 975 ICV_35 $T=28930 1000 0 0 $X=28815 $Y=885
X7773 585 188 VSS VDD 758 188 251 585 ICV_36 $T=16580 43000 0 0 $X=16465 $Y=42885
X7774 53 148 VSS VDD 766 148 257 53 ICV_36 $T=16960 31800 0 0 $X=16845 $Y=31685
X7775 611 250 VSS VDD 778 770 250 761 ICV_36 $T=22280 40200 1 0 $X=22165 $Y=38685
X7776 778 254 VSS VDD 868 604 254 599 ICV_36 $T=22660 34600 1 0 $X=22545 $Y=33085
X7777 610 259 VSS VDD 507 244 259 602 ICV_36 $T=23040 29000 0 0 $X=22925 $Y=28885
X7778 785 268 VSS VDD 786 617 268 612 ICV_36 $T=24560 26200 1 0 $X=24445 $Y=24685
X7779 626 292 VSS VDD 627 292 330 626 ICV_36 $T=26840 9400 0 0 $X=26725 $Y=9285
X7780 629 303 VSS VDD 630 508 303 619 ICV_36 $T=27980 12200 0 0 $X=27865 $Y=12085
X7781 914 739 VDD 738 744 561 VSS ICV_37 $T=9360 43000 0 0 $X=9245 $Y=42885
X7782 736 747 VDD 562 568 564 VSS ICV_37 $T=10880 45800 0 0 $X=10765 $Y=45685
X7783 735 931 VDD 587 590 758 VSS ICV_37 $T=16770 43000 1 0 $X=16655 $Y=41485
X7784 746 757 VDD 759 865 766 VSS ICV_37 $T=18100 34600 1 0 $X=17985 $Y=33085
X7785 734 765 VDD 761 596 770 VSS ICV_37 $T=18480 40200 1 0 $X=18365 $Y=38685
X7786 897 767 VDD 762 222 771 VSS ICV_37 $T=18670 37400 1 0 $X=18555 $Y=35885
X7787 769 593 VDD 592 866 595 VSS ICV_37 $T=19430 37400 0 0 $X=19315 $Y=37285
X7788 764 773 VDD 777 867 780 VSS ICV_37 $T=22470 26200 1 0 $X=22355 $Y=24685
X7789 899 603 VDD 936 616 614 VSS ICV_37 $T=23230 15000 0 0 $X=23115 $Y=14885
X7790 609 933 VDD 612 869 617 VSS ICV_37 $T=23420 23400 0 0 $X=23305 $Y=23285
X7791 779 776 VDD 781 621 784 VSS ICV_37 $T=23610 15000 1 0 $X=23495 $Y=13485
X7792 618 935 VDD 619 954 508 VSS ICV_37 $T=24750 12200 1 0 $X=24635 $Y=10685
X7793 788 937 VDD 789 872 627 VSS ICV_37 $T=26650 9400 1 0 $X=26535 $Y=7885
X7794 77 638 76 VSS VDD 585 76 77 66 ICV_38 $T=5370 43000 0 0 $X=5255 $Y=42885
X7795 78 638 50 VSS VDD 926 50 78 536 ICV_38 $T=5370 45800 1 0 $X=5255 $Y=44285
X7796 84 638 57 VSS VDD 769 57 84 542 ICV_38 $T=5750 37400 1 0 $X=5635 $Y=35885
X7797 110 74 118 VSS VDD 559 97 545 553 ICV_38 $T=8410 12200 1 0 $X=8295 $Y=10685
X7798 161 139 146 VSS VDD 593 146 161 571 ICV_38 $T=13540 37400 1 0 $X=13425 $Y=35885
X7799 201 638 207 VSS VDD 764 207 201 861 ICV_38 $T=17530 26200 1 0 $X=17415 $Y=24685
X7800 220 139 210 VSS VDD 244 210 220 760 ICV_38 $T=19430 29000 1 0 $X=19315 $Y=27485
X7801 229 139 234 VSS VDD 773 234 229 864 ICV_38 $T=20000 26200 1 0 $X=19885 $Y=24685
X7802 237 139 218 VSS VDD 603 218 237 594 ICV_38 $T=20760 15000 0 0 $X=20645 $Y=14885
X7803 274 333 296 VSS VDD 320 274 296 870 ICV_38 $T=26460 31800 0 0 $X=26345 $Y=31685
X7806 VSS VDD b[15] 18 a[15] 43 ICV_39 $T=1950 15000 1 0 $X=1835 $Y=13485
X7807 VSS VDD b[4] 18 a[4] 923 ICV_39 $T=1950 23400 0 0 $X=1835 $Y=23285
X7808 VSS VDD a[11] 37 b[11] 103 ICV_39 $T=1950 29000 0 0 $X=1835 $Y=28885
X7809 VSS VDD a[1] 37 b[1] 56 ICV_39 $T=1950 34600 1 0 $X=1835 $Y=33085
X7810 VSS VDD b[10] 18 a[10] 106 ICV_39 $T=1950 34600 0 0 $X=1835 $Y=34485
X7811 VSS VDD a[9] 37 b[9] 80 ICV_39 $T=1950 37400 0 0 $X=1835 $Y=37285
X7812 VSS VDD a[8] 37 b[8] 76 ICV_39 $T=1950 43000 1 0 $X=1835 $Y=41485
X7813 VSS VDD a[7] 37 b[7] 50 ICV_39 $T=1950 43000 0 0 $X=1835 $Y=42885
X7814 VSS VDD a[6] 37 b[6] 45 ICV_39 $T=1950 45800 1 0 $X=1835 $Y=44285
X7815 VSS VDD 239 638 247 618 ICV_39 $T=21900 3800 0 0 $X=21785 $Y=3685
X7816 VSS VDD 240 139 232 776 ICV_39 $T=21900 15000 1 0 $X=21785 $Y=13485
X7817 VSS VDD 241 139 212 261 ICV_39 $T=21900 17800 0 0 $X=21785 $Y=17685
.ENDS
***************************************
