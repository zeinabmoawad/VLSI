/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sun Dec 11 23:17:47 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 818263663 */

module datapath(in2, in1, out);
   input [31:0]in2;
   input [31:0]in1;
   output [63:0]out;

   HA_X1 i_0 (.A(n_1030), .B(n_1045), .CO(n_1053), .S(n_1052));
   FA_X1 i_1 (.A(n_1040), .B(n_1046), .CI(n_1063), .CO(n_1069), .S(n_1068));
   HA_X1 i_2 (.A(n_1056), .B(n_1053), .CO(n_1071), .S(n_1070));
   HA_X1 i_3 (.A(n_1071), .B(n_1069), .CO(n_1097), .S(n_1096));
   FA_X1 i_5 (.A(n_1107), .B(n_1100), .CI(n_1097), .CO(n_1123), .S(n_1122));
   FA_X1 i_7 (.A(n_1108), .B(n_1101), .CI(n_1114), .CO(n_1148), .S(n_1147));
   FA_X1 i_8 (.A(n_1142), .B(n_1135), .CI(n_1128), .CO(n_1150), .S(n_1149));
   FA_X1 i_9 (.A(n_1147), .B(n_600), .CI(n_603), .CO(n_1152), .S(n_1151));
   HA_X1 i_10 (.A(n_1123), .B(n_1149), .CO(n_1154), .S(n_1153));
   FA_X1 i_11 (.A(n_1129), .B(n_1171), .CI(n_1164), .CO(n_1185), .S(n_1184));
   FA_X1 i_1173 (.A(n_1157), .B(n_1148), .CI(n_572), .CO(n_1187), .S(n_1186));
   FA_X1 i_1174 (.A(n_1150), .B(n_1184), .CI(n_1186), .CO(n_1189), .S(n_1188));
   HA_X1 i_12 (.A(n_1154), .B(n_1152), .CO(n_1191), .S(n_1190));
   FA_X1 i_13 (.A(n_1165), .B(n_1158), .CI(n_1179), .CO(n_1222), .S(n_1221));
   FA_X1 i_14 (.A(n_1214), .B(n_1208), .CI(n_1201), .CO(n_1224), .S(n_1223));
   FA_X1 i_15 (.A(n_1194), .B(n_1221), .CI(n_1185), .CO(n_1226), .S(n_1225));
   FA_X1 i_1208 (.A(n_1187), .B(n_1223), .CI(n_1225), .CO(n_1228), .S(n_1227));
   HA_X1 i_1209 (.A(n_1191), .B(n_1189), .CO(n_1230), .S(n_1229));
   FA_X1 i_16 (.A(n_1209), .B(n_1202), .CI(n_1195), .CO(n_1260), .S(n_1259));
   FA_X1 i_18 (.A(n_1215), .B(n_1254), .CI(n_1247), .CO(n_1262), .S(n_1261));
   FA_X1 i_19 (.A(n_1240), .B(n_1233), .CI(n_1222), .CO(n_1264), .S(n_1263));
   FA_X1 i_20 (.A(n_1259), .B(n_1224), .CI(n_1226), .CO(n_1266), .S(n_1265));
   FA_X1 i_23 (.A(n_1263), .B(n_1261), .CI(n_1265), .CO(n_1268), .S(n_1267));
   HA_X1 i_1243 (.A(n_1230), .B(n_1228), .CO(n_1270), .S(n_1269));
   FA_X1 i_25 (.A(n_1241), .B(n_1234), .CI(n_1260), .CO(n_1308), .S(n_1307));
   FA_X1 i_27 (.A(n_1294), .B(n_1287), .CI(n_1280), .CO(n_1310), .S(n_1309));
   FA_X1 i_28 (.A(n_1273), .B(n_1307), .CI(n_1301), .CO(n_1312), .S(n_1311));
   FA_X1 i_29 (.A(n_1262), .B(n_1264), .CI(n_1309), .CO(n_1314), .S(n_1313));
   FA_X1 i_30 (.A(n_1266), .B(n_1311), .CI(n_1313), .CO(n_1316), .S(n_1315));
   HA_X1 i_1285 (.A(n_1268), .B(n_1270), .CO(n_1318), .S(n_1317));
   FA_X1 i_31 (.A(n_1288), .B(n_1281), .CI(n_1274), .CO(n_1356), .S(n_1355));
   FA_X1 i_32 (.A(n_1302), .B(n_1348), .CI(n_1342), .CO(n_1358), .S(n_1357));
   FA_X1 i_33 (.A(n_1335), .B(n_1328), .CI(n_1321), .CO(n_1360), .S(n_1359));
   FA_X1 i_34 (.A(n_1308), .B(n_1355), .CI(n_1310), .CO(n_1362), .S(n_1361));
   FA_X1 i_35 (.A(n_1312), .B(n_1359), .CI(n_1357), .CO(n_1364), .S(n_1363));
   FA_X1 i_36 (.A(n_1361), .B(n_1314), .CI(n_1316), .CO(n_1366), .S(n_1365));
   HA_X1 i_37 (.A(n_1363), .B(n_1318), .CO(n_1368), .S(n_1367));
   FA_X1 i_38 (.A(n_1343), .B(n_1336), .CI(n_1329), .CO(n_1405), .S(n_1404));
   FA_X1 i_39 (.A(n_1322), .B(n_1356), .CI(n_1349), .CO(n_1407), .S(n_1406));
   FA_X1 i_40 (.A(n_1399), .B(n_1392), .CI(n_1385), .CO(n_1409), .S(n_1408));
   FA_X1 i_41 (.A(n_1378), .B(n_1371), .CI(n_1404), .CO(n_1411), .S(n_1410));
   FA_X1 i_42 (.A(n_1360), .B(n_1358), .CI(n_1406), .CO(n_1413), .S(n_1412));
   FA_X1 i_43 (.A(n_1362), .B(n_1410), .CI(n_1408), .CO(n_1415), .S(n_1414));
   FA_X1 i_44 (.A(n_1412), .B(n_1364), .CI(n_1414), .CO(n_1417), .S(n_1416));
   HA_X1 i_45 (.A(n_1366), .B(n_1368), .CO(n_1419), .S(n_1418));
   FA_X1 i_46 (.A(n_1386), .B(n_1379), .CI(n_1372), .CO(n_1464), .S(n_1463));
   FA_X1 i_47 (.A(n_1405), .B(n_1450), .CI(n_1443), .CO(n_1466), .S(n_1465));
   FA_X1 i_48 (.A(n_1436), .B(n_1429), .CI(n_1422), .CO(n_1468), .S(n_1467));
   FA_X1 i_49 (.A(n_1407), .B(n_1463), .CI(n_1457), .CO(n_1470), .S(n_1469));
   FA_X1 i_50 (.A(n_1409), .B(n_1411), .CI(n_1467), .CO(n_1472), .S(n_1471));
   FA_X1 i_51 (.A(n_1465), .B(n_1413), .CI(n_1469), .CO(n_1474), .S(n_1473));
   FA_X1 i_52 (.A(n_1415), .B(n_1471), .CI(n_1473), .CO(n_1476), .S(n_1475));
   HA_X1 i_53 (.A(n_1417), .B(n_1419), .CO(n_1478), .S(n_1477));
   FA_X1 i_54 (.A(n_1444), .B(n_1437), .CI(n_1430), .CO(n_1523), .S(n_1522));
   FA_X1 i_55 (.A(n_1423), .B(n_1464), .CI(n_1458), .CO(n_1525), .S(n_1524));
   FA_X1 i_56 (.A(n_1515), .B(n_1509), .CI(n_1502), .CO(n_1527), .S(n_1526));
   FA_X1 i_57 (.A(n_1495), .B(n_1488), .CI(n_1481), .CO(n_1529), .S(n_1528));
   FA_X1 i_58 (.A(n_1522), .B(n_1468), .CI(n_1466), .CO(n_1531), .S(n_1530));
   FA_X1 i_59 (.A(n_1524), .B(n_1470), .CI(n_1528), .CO(n_1533), .S(n_1532));
   FA_X1 i_60 (.A(n_1526), .B(n_1530), .CI(n_1472), .CO(n_1535), .S(n_1534));
   FA_X1 i_61 (.A(n_1532), .B(n_1474), .CI(n_1534), .CO(n_1537), .S(n_1536));
   HA_X1 i_62 (.A(n_1476), .B(n_1478), .CO(n_1539), .S(n_1538));
   FA_X1 i_63 (.A(n_1510), .B(n_1503), .CI(n_1496), .CO(n_1583), .S(n_1582));
   FA_X1 i_64 (.A(n_1489), .B(n_1482), .CI(n_1523), .CO(n_1585), .S(n_1584));
   FA_X1 i_65 (.A(n_1516), .B(n_1577), .CI(n_1570), .CO(n_1587), .S(n_1586));
   FA_X1 i_66 (.A(n_1563), .B(n_1556), .CI(n_1549), .CO(n_1589), .S(n_1588));
   FA_X1 i_67 (.A(n_1542), .B(n_1525), .CI(n_1584), .CO(n_1591), .S(n_1590));
   FA_X1 i_68 (.A(n_1582), .B(n_1529), .CI(n_1527), .CO(n_1593), .S(n_1592));
   FA_X1 i_69 (.A(n_1531), .B(n_1588), .CI(n_1586), .CO(n_1595), .S(n_1594));
   FA_X1 i_70 (.A(n_1590), .B(n_1592), .CI(n_1533), .CO(n_1597), .S(n_1596));
   FA_X1 i_71 (.A(n_1535), .B(n_1594), .CI(n_1596), .CO(n_1599), .S(n_1598));
   HA_X1 i_72 (.A(n_1537), .B(n_1539), .CO(n_1601), .S(n_1600));
   FA_X1 i_73 (.A(n_1564), .B(n_1557), .CI(n_1550), .CO(n_1653), .S(n_1652));
   FA_X1 i_74 (.A(n_1543), .B(n_1583), .CI(n_1639), .CO(n_1655), .S(n_1654));
   FA_X1 i_75 (.A(n_1632), .B(n_1625), .CI(n_1618), .CO(n_1657), .S(n_1656));
   FA_X1 i_76 (.A(n_1611), .B(n_1604), .CI(n_1585), .CO(n_1659), .S(n_1658));
   FA_X1 i_77 (.A(n_1652), .B(n_1646), .CI(n_1589), .CO(n_1661), .S(n_1660));
   FA_X1 i_78 (.A(n_1587), .B(n_1654), .CI(n_1593), .CO(n_1663), .S(n_1662));
   FA_X1 i_79 (.A(n_1591), .B(n_1658), .CI(n_1656), .CO(n_1665), .S(n_1664));
   FA_X1 i_80 (.A(n_1660), .B(n_1595), .CI(n_1662), .CO(n_1667), .S(n_1666));
   FA_X1 i_81 (.A(n_1597), .B(n_1664), .CI(n_1666), .CO(n_1669), .S(n_1668));
   HA_X1 i_82 (.A(n_1599), .B(n_1668), .CO(n_1671), .S(n_1670));
   FA_X1 i_83 (.A(n_1633), .B(n_1626), .CI(n_1619), .CO(n_1723), .S(n_1722));
   FA_X1 i_84 (.A(n_1612), .B(n_1605), .CI(n_1653), .CO(n_1725), .S(n_1724));
   FA_X1 i_85 (.A(n_1647), .B(n_1715), .CI(n_1709), .CO(n_1727), .S(n_1726));
   FA_X1 i_86 (.A(n_1702), .B(n_1695), .CI(n_1688), .CO(n_1729), .S(n_1728));
   FA_X1 i_87 (.A(n_1681), .B(n_1674), .CI(n_1724), .CO(n_1731), .S(n_1730));
   FA_X1 i_88 (.A(n_1722), .B(n_1657), .CI(n_1655), .CO(n_1733), .S(n_1732));
   FA_X1 i_89 (.A(n_1659), .B(n_1661), .CI(n_1730), .CO(n_1735), .S(n_1734));
   FA_X1 i_90 (.A(n_1728), .B(n_1726), .CI(n_1663), .CO(n_1737), .S(n_1736));
   FA_X1 i_91 (.A(n_1732), .B(n_1665), .CI(n_1734), .CO(n_1739), .S(n_1738));
   FA_X1 i_92 (.A(n_1736), .B(n_1667), .CI(n_1738), .CO(n_1741), .S(n_1740));
   HA_X1 i_93 (.A(n_1669), .B(n_1740), .CO(n_1743), .S(n_1742));
   FA_X1 i_94 (.A(n_1710), .B(n_1703), .CI(n_1696), .CO(n_1794), .S(n_1793));
   FA_X1 i_95 (.A(n_1689), .B(n_1682), .CI(n_1675), .CO(n_1796), .S(n_1795));
   FA_X1 i_96 (.A(n_1723), .B(n_1716), .CI(n_1788), .CO(n_1798), .S(n_1797));
   FA_X1 i_97 (.A(n_1781), .B(n_1774), .CI(n_1767), .CO(n_1800), .S(n_1799));
   FA_X1 i_98 (.A(n_1760), .B(n_1753), .CI(n_1746), .CO(n_1802), .S(n_1801));
   FA_X1 i_99 (.A(n_1725), .B(n_1795), .CI(n_1793), .CO(n_1804), .S(n_1803));
   FA_X1 i_100 (.A(n_1729), .B(n_1727), .CI(n_1797), .CO(n_1806), .S(n_1805));
   FA_X1 i_101 (.A(n_1733), .B(n_1731), .CI(n_1801), .CO(n_1808), .S(n_1807));
   FA_X1 i_102 (.A(n_1799), .B(n_1805), .CI(n_1803), .CO(n_1810), .S(n_1809));
   FA_X1 i_103 (.A(n_1735), .B(n_1737), .CI(n_1807), .CO(n_1812), .S(n_1811));
   FA_X1 i_104 (.A(n_1739), .B(n_1809), .CI(n_1811), .CO(n_1814), .S(n_1813));
   HA_X1 i_105 (.A(n_1741), .B(n_1743), .CO(n_1816), .S(n_1815));
   FA_X1 i_106 (.A(n_1775), .B(n_1768), .CI(n_1761), .CO(n_1875), .S(n_1874));
   FA_X1 i_107 (.A(n_1754), .B(n_1747), .CI(n_1796), .CO(n_1877), .S(n_1876));
   FA_X1 i_108 (.A(n_1794), .B(n_1861), .CI(n_1854), .CO(n_1879), .S(n_1878));
   FA_X1 i_109 (.A(n_1847), .B(n_1840), .CI(n_1833), .CO(n_1881), .S(n_1880));
   FA_X1 i_110 (.A(n_1826), .B(n_1819), .CI(n_1876), .CO(n_1883), .S(n_1882));
   FA_X1 i_111 (.A(n_1874), .B(n_1868), .CI(n_1802), .CO(n_1885), .S(n_1884));
   FA_X1 i_112 (.A(n_1800), .B(n_1798), .CI(n_1804), .CO(n_1887), .S(n_1886));
   FA_X1 i_113 (.A(n_1882), .B(n_1880), .CI(n_1878), .CO(n_1889), .S(n_1888));
   FA_X1 i_114 (.A(n_1806), .B(n_1886), .CI(n_1884), .CO(n_1891), .S(n_1890));
   FA_X1 i_115 (.A(n_1808), .B(n_1810), .CI(n_1888), .CO(n_1893), .S(n_1892));
   FA_X1 i_116 (.A(n_1812), .B(n_1890), .CI(n_1892), .CO(n_1895), .S(n_1894));
   HA_X1 i_117 (.A(n_1814), .B(n_1894), .CO(n_1897), .S(n_1896));
   FA_X1 i_118 (.A(n_1855), .B(n_1848), .CI(n_1841), .CO(n_1956), .S(n_1955));
   FA_X1 i_119 (.A(n_1834), .B(n_1827), .CI(n_1820), .CO(n_1958), .S(n_1957));
   FA_X1 i_120 (.A(n_1875), .B(n_1869), .CI(n_1948), .CO(n_1960), .S(n_1959));
   FA_X1 i_121 (.A(n_1942), .B(n_1935), .CI(n_1928), .CO(n_1962), .S(n_1961));
   FA_X1 i_122 (.A(n_1921), .B(n_1914), .CI(n_1907), .CO(n_1964), .S(n_1963));
   FA_X1 i_123 (.A(n_1900), .B(n_1877), .CI(n_1957), .CO(n_1966), .S(n_1965));
   FA_X1 i_124 (.A(n_1955), .B(n_1881), .CI(n_1879), .CO(n_1968), .S(n_1967));
   FA_X1 i_125 (.A(n_1959), .B(n_1885), .CI(n_1883), .CO(n_1970), .S(n_1969));
   FA_X1 i_126 (.A(n_1963), .B(n_1961), .CI(n_1965), .CO(n_1972), .S(n_1971));
   FA_X1 i_127 (.A(n_1887), .B(n_1967), .CI(n_1889), .CO(n_1974), .S(n_1973));
   FA_X1 i_128 (.A(n_1969), .B(n_1891), .CI(n_1971), .CO(n_1976), .S(n_1975));
   FA_X1 i_129 (.A(n_1973), .B(n_1893), .CI(n_1975), .CO(n_1978), .S(n_1977));
   HA_X1 i_130 (.A(n_1895), .B(n_1977), .CO(n_1980), .S(n_1979));
   FA_X1 i_131 (.A(n_1943), .B(n_1936), .CI(n_1929), .CO(n_2038), .S(n_2037));
   FA_X1 i_132 (.A(n_1922), .B(n_1915), .CI(n_1908), .CO(n_2040), .S(n_2039));
   FA_X1 i_133 (.A(n_1901), .B(n_1958), .CI(n_1956), .CO(n_2042), .S(n_2041));
   FA_X1 i_134 (.A(n_1949), .B(n_2032), .CI(n_2025), .CO(n_2044), .S(n_2043));
   FA_X1 i_135 (.A(n_2018), .B(n_2011), .CI(n_2004), .CO(n_2046), .S(n_2045));
   FA_X1 i_136 (.A(n_1997), .B(n_1990), .CI(n_1983), .CO(n_2048), .S(n_2047));
   FA_X1 i_137 (.A(n_2039), .B(n_2037), .CI(n_1964), .CO(n_2050), .S(n_2049));
   FA_X1 i_138 (.A(n_1962), .B(n_1960), .CI(n_2041), .CO(n_2052), .S(n_2051));
   FA_X1 i_139 (.A(n_1968), .B(n_1966), .CI(n_2047), .CO(n_2054), .S(n_2053));
   FA_X1 i_140 (.A(n_2045), .B(n_2043), .CI(n_1970), .CO(n_2056), .S(n_2055));
   FA_X1 i_141 (.A(n_2051), .B(n_2049), .CI(n_1972), .CO(n_2058), .S(n_2057));
   FA_X1 i_142 (.A(n_2053), .B(n_1974), .CI(n_2055), .CO(n_2060), .S(n_2059));
   FA_X1 i_143 (.A(n_2057), .B(n_1976), .CI(n_2059), .CO(n_2062), .S(n_2061));
   HA_X1 i_144 (.A(n_1978), .B(n_2061), .CO(n_2064), .S(n_2063));
   FA_X1 i_145 (.A(n_2019), .B(n_2012), .CI(n_2005), .CO(n_2130), .S(n_2129));
   FA_X1 i_146 (.A(n_1998), .B(n_1991), .CI(n_1984), .CO(n_2132), .S(n_2131));
   FA_X1 i_147 (.A(n_2040), .B(n_2038), .CI(n_2116), .CO(n_2134), .S(n_2133));
   FA_X1 i_148 (.A(n_2109), .B(n_2102), .CI(n_2095), .CO(n_2136), .S(n_2135));
   FA_X1 i_149 (.A(n_2088), .B(n_2081), .CI(n_2074), .CO(n_2138), .S(n_2137));
   FA_X1 i_150 (.A(n_2067), .B(n_2042), .CI(n_2131), .CO(n_2140), .S(n_2139));
   FA_X1 i_151 (.A(n_2129), .B(n_2123), .CI(n_2048), .CO(n_2142), .S(n_2141));
   FA_X1 i_152 (.A(n_2046), .B(n_2044), .CI(n_2133), .CO(n_2144), .S(n_2143));
   FA_X1 i_153 (.A(n_2050), .B(n_2137), .CI(n_2135), .CO(n_2146), .S(n_2145));
   FA_X1 i_154 (.A(n_2139), .B(n_2052), .CI(n_2143), .CO(n_2148), .S(n_2147));
   FA_X1 i_155 (.A(n_2141), .B(n_2054), .CI(n_2056), .CO(n_2150), .S(n_2149));
   FA_X1 i_156 (.A(n_2058), .B(n_2145), .CI(n_2147), .CO(n_2152), .S(n_2151));
   FA_X1 i_157 (.A(n_2149), .B(n_2060), .CI(n_2151), .CO(n_2154), .S(n_2153));
   HA_X1 i_158 (.A(n_2062), .B(n_2153), .CO(n_2156), .S(n_2155));
   FA_X1 i_159 (.A(n_2110), .B(n_2103), .CI(n_2096), .CO(n_2222), .S(n_2221));
   FA_X1 i_160 (.A(n_2089), .B(n_2082), .CI(n_2075), .CO(n_2224), .S(n_2223));
   FA_X1 i_161 (.A(n_2068), .B(n_2132), .CI(n_2130), .CO(n_2226), .S(n_2225));
   FA_X1 i_162 (.A(n_2124), .B(n_2214), .CI(n_2208), .CO(n_2228), .S(n_2227));
   FA_X1 i_163 (.A(n_2201), .B(n_2194), .CI(n_2187), .CO(n_2230), .S(n_2229));
   FA_X1 i_164 (.A(n_2180), .B(n_2173), .CI(n_2166), .CO(n_2232), .S(n_2231));
   FA_X1 i_165 (.A(n_2159), .B(n_2223), .CI(n_2221), .CO(n_2234), .S(n_2233));
   FA_X1 i_166 (.A(n_2138), .B(n_2136), .CI(n_2134), .CO(n_2236), .S(n_2235));
   FA_X1 i_167 (.A(n_2225), .B(n_2142), .CI(n_2140), .CO(n_2238), .S(n_2237));
   FA_X1 i_168 (.A(n_2231), .B(n_2229), .CI(n_2227), .CO(n_2240), .S(n_2239));
   FA_X1 i_169 (.A(n_2144), .B(n_2235), .CI(n_2233), .CO(n_2242), .S(n_2241));
   FA_X1 i_170 (.A(n_2146), .B(n_2237), .CI(n_2148), .CO(n_2244), .S(n_2243));
   FA_X1 i_171 (.A(n_2150), .B(n_2239), .CI(n_2241), .CO(n_2246), .S(n_2245));
   FA_X1 i_172 (.A(n_2152), .B(n_2243), .CI(n_2245), .CO(n_2248), .S(n_2247));
   HA_X1 i_173 (.A(n_2154), .B(n_2156), .CO(n_2250), .S(n_2249));
   FA_X1 i_174 (.A(n_2209), .B(n_2202), .CI(n_2195), .CO(n_2315), .S(n_2314));
   FA_X1 i_175 (.A(n_2188), .B(n_2181), .CI(n_2174), .CO(n_2317), .S(n_2316));
   FA_X1 i_176 (.A(n_2167), .B(n_2160), .CI(n_2224), .CO(n_2319), .S(n_2318));
   FA_X1 i_177 (.A(n_2222), .B(n_2215), .CI(n_2309), .CO(n_2321), .S(n_2320));
   FA_X1 i_178 (.A(n_2302), .B(n_2295), .CI(n_2288), .CO(n_2323), .S(n_2322));
   FA_X1 i_179 (.A(n_2281), .B(n_2274), .CI(n_2267), .CO(n_2325), .S(n_2324));
   FA_X1 i_180 (.A(n_2260), .B(n_2253), .CI(n_2226), .CO(n_2327), .S(n_2326));
   FA_X1 i_181 (.A(n_2318), .B(n_2316), .CI(n_2314), .CO(n_2329), .S(n_2328));
   FA_X1 i_182 (.A(n_2232), .B(n_2230), .CI(n_2228), .CO(n_2331), .S(n_2330));
   FA_X1 i_183 (.A(n_2320), .B(n_2236), .CI(n_2234), .CO(n_2333), .S(n_2332));
   FA_X1 i_184 (.A(n_2326), .B(n_2324), .CI(n_2322), .CO(n_2335), .S(n_2334));
   FA_X1 i_185 (.A(n_2238), .B(n_2330), .CI(n_2328), .CO(n_2337), .S(n_2336));
   FA_X1 i_186 (.A(n_2240), .B(n_2332), .CI(n_2242), .CO(n_2339), .S(n_2338));
   FA_X1 i_187 (.A(n_2334), .B(n_2244), .CI(n_2336), .CO(n_2341), .S(n_2340));
   FA_X1 i_188 (.A(n_2338), .B(n_2246), .CI(n_2340), .CO(n_2343), .S(n_2342));
   HA_X1 i_189 (.A(n_2248), .B(n_2342), .CO(n_2345), .S(n_2344));
   FA_X1 i_190 (.A(n_2296), .B(n_2289), .CI(n_2282), .CO(n_2418), .S(n_2417));
   FA_X1 i_191 (.A(n_2275), .B(n_2268), .CI(n_2261), .CO(n_2420), .S(n_2419));
   FA_X1 i_192 (.A(n_2254), .B(n_2317), .CI(n_2315), .CO(n_2422), .S(n_2421));
   FA_X1 i_193 (.A(n_2404), .B(n_2397), .CI(n_2390), .CO(n_2424), .S(n_2423));
   FA_X1 i_194 (.A(n_2383), .B(n_2376), .CI(n_2369), .CO(n_2426), .S(n_2425));
   FA_X1 i_195 (.A(n_2362), .B(n_2355), .CI(n_2348), .CO(n_2428), .S(n_2427));
   FA_X1 i_196 (.A(n_2319), .B(n_2419), .CI(n_2417), .CO(n_2430), .S(n_2429));
   FA_X1 i_197 (.A(n_2411), .B(n_2325), .CI(n_2323), .CO(n_2432), .S(n_2431));
   FA_X1 i_198 (.A(n_2321), .B(n_2327), .CI(n_2421), .CO(n_2434), .S(n_2433));
   FA_X1 i_199 (.A(n_2331), .B(n_2329), .CI(n_2427), .CO(n_2436), .S(n_2435));
   FA_X1 i_200 (.A(n_2425), .B(n_2423), .CI(n_2333), .CO(n_2438), .S(n_2437));
   FA_X1 i_201 (.A(n_2431), .B(n_2429), .CI(n_2335), .CO(n_2440), .S(n_2439));
   FA_X1 i_202 (.A(n_2433), .B(n_2435), .CI(n_2337), .CO(n_2442), .S(n_2441));
   FA_X1 i_203 (.A(n_2437), .B(n_2339), .CI(n_2439), .CO(n_2444), .S(n_2443));
   FA_X1 i_204 (.A(n_2441), .B(n_2341), .CI(n_2443), .CO(n_2446), .S(n_2445));
   HA_X1 i_205 (.A(n_2343), .B(n_2445), .CO(n_2448), .S(n_2447));
   FA_X1 i_206 (.A(n_2398), .B(n_2391), .CI(n_2384), .CO(n_2521), .S(n_2520));
   FA_X1 i_207 (.A(n_2377), .B(n_2370), .CI(n_2363), .CO(n_2523), .S(n_2522));
   FA_X1 i_208 (.A(n_2356), .B(n_2349), .CI(n_2420), .CO(n_2525), .S(n_2524));
   FA_X1 i_209 (.A(n_2418), .B(n_2412), .CI(n_2513), .CO(n_2527), .S(n_2526));
   FA_X1 i_210 (.A(n_2507), .B(n_2500), .CI(n_2493), .CO(n_2529), .S(n_2528));
   FA_X1 i_211 (.A(n_2486), .B(n_2479), .CI(n_2472), .CO(n_2531), .S(n_2530));
   FA_X1 i_212 (.A(n_2465), .B(n_2458), .CI(n_2451), .CO(n_2533), .S(n_2532));
   FA_X1 i_213 (.A(n_2422), .B(n_2524), .CI(n_2522), .CO(n_2535), .S(n_2534));
   FA_X1 i_214 (.A(n_2520), .B(n_2428), .CI(n_2426), .CO(n_2537), .S(n_2536));
   FA_X1 i_215 (.A(n_2424), .B(n_2526), .CI(n_2432), .CO(n_2539), .S(n_2538));
   FA_X1 i_216 (.A(n_2430), .B(n_2532), .CI(n_2530), .CO(n_2541), .S(n_2540));
   FA_X1 i_217 (.A(n_2528), .B(n_2434), .CI(n_2536), .CO(n_2543), .S(n_2542));
   FA_X1 i_218 (.A(n_2534), .B(n_2436), .CI(n_2438), .CO(n_2545), .S(n_2544));
   FA_X1 i_219 (.A(n_2538), .B(n_2440), .CI(n_2540), .CO(n_2547), .S(n_2546));
   FA_X1 i_220 (.A(n_2542), .B(n_2442), .CI(n_2544), .CO(n_2549), .S(n_2548));
   FA_X1 i_221 (.A(n_2546), .B(n_2444), .CI(n_2548), .CO(n_2551), .S(n_2550));
   HA_X1 i_222 (.A(n_2446), .B(n_2550), .CO(n_2553), .S(n_2552));
   FA_X1 i_223 (.A(n_2508), .B(n_2501), .CI(n_2494), .CO(n_2625), .S(n_2624));
   FA_X1 i_224 (.A(n_2487), .B(n_2480), .CI(n_2473), .CO(n_2627), .S(n_2626));
   FA_X1 i_225 (.A(n_2466), .B(n_2459), .CI(n_2452), .CO(n_2629), .S(n_2628));
   FA_X1 i_226 (.A(n_2523), .B(n_2521), .CI(n_2514), .CO(n_2631), .S(n_2630));
   FA_X1 i_227 (.A(n_2619), .B(n_2612), .CI(n_2605), .CO(n_2633), .S(n_2632));
   FA_X1 i_228 (.A(n_2598), .B(n_2591), .CI(n_2584), .CO(n_2635), .S(n_2634));
   FA_X1 i_229 (.A(n_2577), .B(n_2570), .CI(n_2563), .CO(n_2637), .S(n_2636));
   FA_X1 i_230 (.A(n_2556), .B(n_2525), .CI(n_2628), .CO(n_2639), .S(n_2638));
   FA_X1 i_231 (.A(n_2626), .B(n_2624), .CI(n_2533), .CO(n_2641), .S(n_2640));
   FA_X1 i_232 (.A(n_2531), .B(n_2529), .CI(n_2527), .CO(n_2643), .S(n_2642));
   FA_X1 i_233 (.A(n_2630), .B(n_2537), .CI(n_2535), .CO(n_2645), .S(n_2644));
   FA_X1 i_234 (.A(n_2636), .B(n_2634), .CI(n_2632), .CO(n_2647), .S(n_2646));
   FA_X1 i_235 (.A(n_2638), .B(n_2539), .CI(n_2642), .CO(n_2649), .S(n_2648));
   FA_X1 i_236 (.A(n_2640), .B(n_2541), .CI(n_2644), .CO(n_2651), .S(n_2650));
   FA_X1 i_237 (.A(n_2543), .B(n_2545), .CI(n_2646), .CO(n_2653), .S(n_2652));
   FA_X1 i_238 (.A(n_2648), .B(n_2650), .CI(n_2547), .CO(n_2655), .S(n_2654));
   FA_X1 i_239 (.A(n_2549), .B(n_2652), .CI(n_2654), .CO(n_2657), .S(n_2656));
   HA_X1 i_240 (.A(n_2551), .B(n_2656), .CO(n_2659), .S(n_2658));
   FA_X1 i_241 (.A(n_2564), .B(n_2557), .CI(n_2629), .CO(n_2743), .S(n_2742));
   FA_X1 i_242 (.A(n_2627), .B(n_2625), .CI(n_2725), .CO(n_2745), .S(n_2744));
   FA_X1 i_243 (.A(n_2718), .B(n_2711), .CI(n_2704), .CO(n_2747), .S(n_2746));
   FA_X1 i_244 (.A(n_2697), .B(n_2690), .CI(n_2683), .CO(n_2749), .S(n_2748));
   FA_X1 i_245 (.A(n_2676), .B(n_2669), .CI(n_2662), .CO(n_2751), .S(n_2750));
   FA_X1 i_246 (.A(n_2631), .B(n_2742), .CI(n_1442), .CO(n_2753), .S(n_2752));
   FA_X1 i_247 (.A(n_1445), .B(n_2732), .CI(n_2637), .CO(n_2755), .S(n_2754));
   FA_X1 i_248 (.A(n_2635), .B(n_2633), .CI(n_2744), .CO(n_2757), .S(n_2756));
   FA_X1 i_249 (.A(n_2643), .B(n_2641), .CI(n_2639), .CO(n_2759), .S(n_2758));
   FA_X1 i_250 (.A(n_2750), .B(n_2748), .CI(n_2746), .CO(n_2761), .S(n_2760));
   FA_X1 i_251 (.A(n_2645), .B(n_2756), .CI(n_2754), .CO(n_2763), .S(n_2762));
   FA_X1 i_252 (.A(n_2752), .B(n_2647), .CI(n_2758), .CO(n_2765), .S(n_2764));
   FA_X1 i_253 (.A(n_2649), .B(n_2760), .CI(n_2651), .CO(n_2767), .S(n_2766));
   FA_X1 i_254 (.A(n_2764), .B(n_2762), .CI(n_2653), .CO(n_2769), .S(n_2768));
   FA_X1 i_255 (.A(n_2655), .B(n_2766), .CI(n_2768), .CO(n_2771), .S(n_2770));
   HA_X1 i_256 (.A(n_2657), .B(n_2770), .CO(n_2773), .S(n_2772));
   FA_X1 i_257 (.A(n_2847), .B(n_2840), .CI(n_2833), .CO(n_2862), .S(n_2861));
   FA_X1 i_258 (.A(n_2784), .B(n_2775), .CI(n_2743), .CO(n_2868), .S(n_2867));
   FA_X1 i_259 (.A(n_1691), .B(n_1692), .CI(n_1693), .CO(n_2870), .S(n_2869));
   FA_X1 i_260 (.A(n_2751), .B(n_2749), .CI(n_2747), .CO(n_2872), .S(n_2871));
   FA_X1 i_261 (.A(n_2745), .B(n_1446), .CI(n_2755), .CO(n_2874), .S(n_2873));
   FA_X1 i_262 (.A(n_2753), .B(n_2867), .CI(n_1439), .CO(n_2876), .S(n_2875));
   FA_X1 i_263 (.A(n_1440), .B(n_2861), .CI(n_2759), .CO(n_2878), .S(n_2877));
   FA_X1 i_264 (.A(n_2757), .B(n_2871), .CI(n_2869), .CO(n_2880), .S(n_2879));
   FA_X1 i_265 (.A(n_2761), .B(n_2873), .CI(n_2763), .CO(n_2882), .S(n_2881));
   FA_X1 i_266 (.A(n_2877), .B(n_2875), .CI(n_2765), .CO(n_2884), .S(n_2883));
   FA_X1 i_267 (.A(n_2879), .B(n_2767), .CI(n_2881), .CO(n_2886), .S(n_2885));
   FA_X1 i_268 (.A(n_2769), .B(n_2883), .CI(n_2885), .CO(n_2888), .S(n_2887));
   HA_X1 i_269 (.A(n_2771), .B(n_2887), .CO(n_2890), .S(n_2889));
   FA_X1 i_270 (.A(n_2848), .B(n_2960), .CI(n_2953), .CO(n_2975), .S(n_2974));
   FA_X1 i_271 (.A(n_2946), .B(n_2939), .CI(n_2932), .CO(n_2977), .S(n_2976));
   FA_X1 i_272 (.A(n_2862), .B(n_2868), .CI(n_1694), .CO(n_2987), .S(n_2986));
   FA_X1 i_273 (.A(n_2872), .B(n_2870), .CI(n_1686), .CO(n_2989), .S(n_2988));
   FA_X1 i_274 (.A(n_1687), .B(n_2976), .CI(n_2974), .CO(n_2991), .S(n_2990));
   FA_X1 i_275 (.A(n_2874), .B(n_1441), .CI(n_1447), .CO(n_2993), .S(n_2992));
   FA_X1 i_276 (.A(n_2876), .B(n_2986), .CI(n_2878), .CO(n_2995), .S(n_2994));
   FA_X1 i_277 (.A(n_2988), .B(n_2880), .CI(n_2990), .CO(n_2997), .S(n_2996));
   FA_X1 i_278 (.A(n_2882), .B(n_2992), .CI(n_2994), .CO(n_2999), .S(n_2998));
   FA_X1 i_279 (.A(n_2884), .B(n_2996), .CI(n_2886), .CO(n_3001), .S(n_3000));
   FA_X1 i_280 (.A(n_2998), .B(n_3000), .CI(n_2888), .CO(n_3003), .S(n_3002));
   FA_X1 i_281 (.A(n_2977), .B(n_2975), .CI(n_715), .CO(n_3097), .S(n_3096));
   FA_X1 i_282 (.A(n_2987), .B(n_3096), .CI(n_1690), .CO(n_3103), .S(n_3102));
   FA_X1 i_283 (.A(n_1697), .B(n_2991), .CI(n_2989), .CO(n_3105), .S(n_3104));
   FA_X1 i_284 (.A(n_1448), .B(n_2993), .CI(n_2995), .CO(n_3107), .S(n_3106));
   FA_X1 i_285 (.A(n_883), .B(n_3104), .CI(n_3102), .CO(n_3109), .S(n_3108));
   FA_X1 i_286 (.A(n_2997), .B(n_3106), .CI(n_2999), .CO(n_3111), .S(n_3110));
   FA_X1 i_287 (.A(n_3108), .B(n_3001), .CI(n_3110), .CO(n_3113), .S(n_3112));
   FA_X1 i_288 (.A(n_3115), .B(n_1387), .CI(n_1832), .CO(n_3201), .S(n_3200));
   FA_X1 i_289 (.A(n_3200), .B(n_1449), .CI(n_3097), .CO(n_3211), .S(n_3210));
   FA_X1 i_290 (.A(n_1698), .B(n_3105), .CI(n_3103), .CO(n_3215), .S(n_3214));
   FA_X1 i_291 (.A(n_1610), .B(n_3210), .CI(n_3107), .CO(n_3217), .S(n_3216));
   FA_X1 i_292 (.A(n_884), .B(n_3214), .CI(n_3109), .CO(n_3219), .S(n_3218));
   FA_X1 i_293 (.A(n_3216), .B(n_3111), .CI(n_3218), .CO(n_3221), .S(n_3220));
   FA_X1 i_294 (.A(n_718), .B(n_3181), .CI(n_3281), .CO(n_3295), .S(n_3294));
   FA_X1 i_295 (.A(n_3274), .B(n_3267), .CI(n_3260), .CO(n_3297), .S(n_3296));
   FA_X1 i_296 (.A(n_3253), .B(n_3246), .CI(n_3239), .CO(n_3299), .S(n_3298));
   FA_X1 i_297 (.A(n_3232), .B(n_3223), .CI(n_1685), .CO(n_3301), .S(n_3300));
   FA_X1 i_298 (.A(n_3294), .B(n_1835), .CI(n_716), .CO(n_3307), .S(n_3306));
   FA_X1 i_299 (.A(n_882), .B(n_3201), .CI(n_3300), .CO(n_3309), .S(n_3308));
   FA_X1 i_300 (.A(n_3298), .B(n_3296), .CI(n_1699), .CO(n_3311), .S(n_3310));
   FA_X1 i_301 (.A(n_3211), .B(n_3308), .CI(n_3306), .CO(n_3315), .S(n_3314));
   FA_X1 i_302 (.A(n_885), .B(n_3310), .CI(n_3215), .CO(n_3317), .S(n_3316));
   FA_X1 i_303 (.A(n_1613), .B(n_3217), .CI(n_3314), .CO(n_3319), .S(n_3318));
   FA_X1 i_304 (.A(n_3316), .B(n_3219), .CI(n_3318), .CO(n_3321), .S(n_3320));
   FA_X1 i_305 (.A(n_3282), .B(n_3275), .CI(n_3268), .CO(n_3388), .S(n_3387));
   FA_X1 i_306 (.A(n_1606), .B(n_1607), .CI(n_1608), .CO(n_3394), .S(n_3393));
   FA_X1 i_307 (.A(n_3380), .B(n_3374), .CI(n_3367), .CO(n_3396), .S(n_3395));
   FA_X1 i_308 (.A(n_3360), .B(n_3353), .CI(n_3346), .CO(n_3398), .S(n_3397));
   FA_X1 i_309 (.A(n_3339), .B(n_3332), .CI(n_3323), .CO(n_3400), .S(n_3399));
   FA_X1 i_310 (.A(n_3387), .B(n_3299), .CI(n_3297), .CO(n_3404), .S(n_3403));
   FA_X1 i_311 (.A(n_3295), .B(n_3301), .CI(n_3393), .CO(n_3406), .S(n_3405));
   FA_X1 i_312 (.A(n_1603), .B(n_1609), .CI(n_3399), .CO(n_3408), .S(n_3407));
   FA_X1 i_313 (.A(n_3397), .B(n_3395), .CI(n_3307), .CO(n_3410), .S(n_3409));
   FA_X1 i_314 (.A(n_3403), .B(n_1838), .CI(n_3309), .CO(n_3412), .S(n_3411));
   FA_X1 i_315 (.A(n_3405), .B(n_3311), .CI(n_3407), .CO(n_3414), .S(n_3413));
   FA_X1 i_316 (.A(n_1614), .B(n_3409), .CI(n_3315), .CO(n_3416), .S(n_3415));
   FA_X1 i_317 (.A(n_3411), .B(n_3413), .CI(n_3317), .CO(n_3418), .S(n_3417));
   FA_X1 i_318 (.A(n_3415), .B(n_3319), .CI(n_3417), .CO(n_3420), .S(n_3419));
   FA_X1 i_319 (.A(n_3333), .B(n_3324), .CI(n_1836), .CO(n_3491), .S(n_3490));
   FA_X1 i_320 (.A(n_1837), .B(n_3388), .CI(n_3480), .CO(n_3493), .S(n_3492));
   FA_X1 i_321 (.A(n_3473), .B(n_3466), .CI(n_3459), .CO(n_3495), .S(n_3494));
   FA_X1 i_322 (.A(n_3452), .B(n_3445), .CI(n_3438), .CO(n_3497), .S(n_3496));
   FA_X1 i_323 (.A(n_3431), .B(n_3422), .CI(n_3394), .CO(n_3499), .S(n_3498));
   FA_X1 i_324 (.A(n_3490), .B(n_1906), .CI(n_1909), .CO(n_3501), .S(n_3500));
   FA_X1 i_325 (.A(n_3400), .B(n_3398), .CI(n_3396), .CO(n_3503), .S(n_3502));
   FA_X1 i_326 (.A(n_3492), .B(n_3404), .CI(n_1839), .CO(n_3505), .S(n_3504));
   FA_X1 i_327 (.A(n_3498), .B(n_3496), .CI(n_3494), .CO(n_3507), .S(n_3506));
   FA_X1 i_328 (.A(n_3406), .B(n_3502), .CI(n_3500), .CO(n_3509), .S(n_3508));
   FA_X1 i_329 (.A(n_3408), .B(n_3410), .CI(n_3504), .CO(n_3511), .S(n_3510));
   FA_X1 i_330 (.A(n_3412), .B(n_3506), .CI(n_3414), .CO(n_3513), .S(n_3512));
   FA_X1 i_331 (.A(n_3508), .B(n_3510), .CI(n_3416), .CO(n_3515), .S(n_3514));
   FA_X1 i_332 (.A(n_3418), .B(n_3512), .CI(n_3514), .CO(n_3517), .S(n_3516));
   FA_X1 i_333 (.A(n_516), .B(n_3474), .CI(n_3467), .CO(n_3576), .S(n_3575));
   FA_X1 i_334 (.A(n_3460), .B(n_3453), .CI(n_3446), .CO(n_3578), .S(n_3577));
   FA_X1 i_335 (.A(n_3570), .B(n_3563), .CI(n_3556), .CO(n_3584), .S(n_3583));
   FA_X1 i_336 (.A(n_3549), .B(n_3542), .CI(n_3535), .CO(n_3586), .S(n_3585));
   FA_X1 i_337 (.A(n_3528), .B(n_3519), .CI(n_3491), .CO(n_3588), .S(n_3587));
   FA_X1 i_338 (.A(n_1911), .B(n_3577), .CI(n_3575), .CO(n_3590), .S(n_3589));
   FA_X1 i_339 (.A(n_3497), .B(n_3495), .CI(n_3493), .CO(n_3592), .S(n_3591));
   FA_X1 i_340 (.A(n_3499), .B(n_1910), .CI(n_3503), .CO(n_3594), .S(n_3593));
   FA_X1 i_341 (.A(n_3501), .B(n_3587), .CI(n_3585), .CO(n_3596), .S(n_3595));
   FA_X1 i_342 (.A(n_3583), .B(n_3505), .CI(n_3591), .CO(n_3598), .S(n_3597));
   FA_X1 i_343 (.A(n_3589), .B(n_3507), .CI(n_3593), .CO(n_3600), .S(n_3599));
   FA_X1 i_344 (.A(n_3509), .B(n_3595), .CI(n_3597), .CO(n_3602), .S(n_3601));
   FA_X1 i_345 (.A(n_3511), .B(n_3599), .CI(n_3513), .CO(n_3604), .S(n_3603));
   FA_X1 i_346 (.A(n_3515), .B(n_3601), .CI(n_3603), .CO(n_3606), .S(n_3605));
   FA_X1 i_347 (.A(n_3571), .B(n_3564), .CI(n_3557), .CO(n_3666), .S(n_3665));
   FA_X1 i_348 (.A(n_3550), .B(n_3543), .CI(n_3536), .CO(n_3668), .S(n_3667));
   FA_X1 i_349 (.A(n_3578), .B(n_3576), .CI(n_3658), .CO(n_3672), .S(n_3671));
   FA_X1 i_350 (.A(n_3652), .B(n_3645), .CI(n_3638), .CO(n_3674), .S(n_3673));
   FA_X1 i_351 (.A(n_3631), .B(n_3624), .CI(n_3617), .CO(n_3676), .S(n_3675));
   FA_X1 i_352 (.A(n_3667), .B(n_3665), .CI(n_3586), .CO(n_3680), .S(n_3679));
   FA_X1 i_353 (.A(n_3584), .B(n_3588), .CI(n_3671), .CO(n_3682), .S(n_3681));
   FA_X1 i_354 (.A(n_3592), .B(n_3590), .CI(n_3675), .CO(n_3684), .S(n_3683));
   FA_X1 i_355 (.A(n_3673), .B(n_1913), .CI(n_3594), .CO(n_3686), .S(n_3685));
   FA_X1 i_356 (.A(n_3679), .B(n_3596), .CI(n_3681), .CO(n_3688), .S(n_3687));
   FA_X1 i_357 (.A(n_3683), .B(n_3598), .CI(n_3685), .CO(n_3690), .S(n_3689));
   FA_X1 i_358 (.A(n_3600), .B(n_3687), .CI(n_3602), .CO(n_3692), .S(n_3691));
   FA_X1 i_359 (.A(n_3689), .B(n_3604), .CI(n_3691), .CO(n_3694), .S(n_3693));
   FA_X1 i_360 (.A(n_3653), .B(n_3646), .CI(n_3639), .CO(n_1), .S(n_0));
   FA_X1 i_361 (.A(n_3632), .B(n_3625), .CI(n_3618), .CO(n_3), .S(n_2));
   FA_X1 i_362 (.A(n_3609), .B(n_3668), .CI(n_3666), .CO(n_5), .S(n_4));
   FA_X1 i_363 (.A(n_398), .B(n_397), .CI(n_3733), .CO(n_7), .S(n_6));
   FA_X1 i_364 (.A(n_3726), .B(n_3719), .CI(n_3712), .CO(n_9), .S(n_8));
   FA_X1 i_365 (.A(n_3705), .B(n_3696), .CI(n_1912), .CO(n_11), .S(n_10));
   FA_X1 i_366 (.A(n_2), .B(n_0), .CI(n_3676), .CO(n_13), .S(n_12));
   FA_X1 i_367 (.A(n_3674), .B(n_3672), .CI(n_4), .CO(n_15), .S(n_14));
   FA_X1 i_368 (.A(n_3680), .B(n_1916), .CI(n_10), .CO(n_17), .S(n_16));
   FA_X1 i_369 (.A(n_8), .B(n_6), .CI(n_3682), .CO(n_19), .S(n_18));
   FA_X1 i_370 (.A(n_14), .B(n_12), .CI(n_3684), .CO(n_21), .S(n_20));
   FA_X1 i_371 (.A(n_3686), .B(n_16), .CI(n_3688), .CO(n_23), .S(n_22));
   FA_X1 i_372 (.A(n_18), .B(n_20), .CI(n_3690), .CO(n_25), .S(n_24));
   FA_X1 i_373 (.A(n_22), .B(n_3692), .CI(n_24), .CO(n_27), .S(n_26));
   FA_X1 i_374 (.A(n_515), .B(n_396), .CI(n_3734), .CO(n_29), .S(n_28));
   FA_X1 i_375 (.A(n_3727), .B(n_3720), .CI(n_3713), .CO(n_31), .S(n_30));
   FA_X1 i_376 (.A(n_3706), .B(n_3697), .CI(n_3), .CO(n_33), .S(n_32));
   FA_X1 i_377 (.A(n_1), .B(n_395), .CI(n_514), .CO(n_35), .S(n_34));
   FA_X1 i_378 (.A(n_513), .B(n_512), .CI(n_511), .CO(n_37), .S(n_36));
   FA_X1 i_379 (.A(n_510), .B(n_509), .CI(n_394), .CO(n_39), .S(n_38));
   FA_X1 i_380 (.A(n_5), .B(n_32), .CI(n_30), .CO(n_41), .S(n_40));
   FA_X1 i_381 (.A(n_28), .B(n_9), .CI(n_7), .CO(n_43), .S(n_42));
   FA_X1 i_382 (.A(n_11), .B(n_34), .CI(n_13), .CO(n_45), .S(n_44));
   FA_X1 i_383 (.A(n_38), .B(n_36), .CI(n_15), .CO(n_47), .S(n_46));
   FA_X1 i_384 (.A(n_42), .B(n_40), .CI(n_17), .CO(n_49), .S(n_48));
   FA_X1 i_385 (.A(n_19), .B(n_44), .CI(n_21), .CO(n_51), .S(n_50));
   FA_X1 i_386 (.A(n_46), .B(n_23), .CI(n_48), .CO(n_53), .S(n_52));
   FA_X1 i_387 (.A(n_50), .B(n_25), .CI(n_52), .CO(n_55), .S(n_54));
   FA_X1 i_388 (.A(n_508), .B(n_507), .CI(n_506), .CO(n_57), .S(n_56));
   FA_X1 i_389 (.A(n_505), .B(n_504), .CI(n_503), .CO(n_59), .S(n_58));
   FA_X1 i_390 (.A(n_391), .B(n_31), .CI(n_29), .CO(n_61), .S(n_60));
   FA_X1 i_391 (.A(n_502), .B(n_501), .CI(n_500), .CO(n_63), .S(n_62));
   FA_X1 i_392 (.A(n_499), .B(n_498), .CI(n_497), .CO(n_65), .S(n_64));
   FA_X1 i_393 (.A(n_496), .B(n_33), .CI(n_58), .CO(n_67), .S(n_66));
   FA_X1 i_394 (.A(n_56), .B(n_39), .CI(n_37), .CO(n_69), .S(n_68));
   FA_X1 i_395 (.A(n_35), .B(n_60), .CI(n_43), .CO(n_71), .S(n_70));
   FA_X1 i_396 (.A(n_41), .B(n_64), .CI(n_62), .CO(n_73), .S(n_72));
   FA_X1 i_397 (.A(n_66), .B(n_45), .CI(n_68), .CO(n_75), .S(n_74));
   FA_X1 i_398 (.A(n_47), .B(n_70), .CI(n_49), .CO(n_77), .S(n_76));
   FA_X1 i_399 (.A(n_72), .B(n_74), .CI(n_51), .CO(n_79), .S(n_78));
   FA_X1 i_400 (.A(n_76), .B(n_53), .CI(n_78), .CO(n_81), .S(n_80));
   FA_X1 i_401 (.A(n_495), .B(n_494), .CI(n_493), .CO(n_83), .S(n_82));
   FA_X1 i_402 (.A(n_492), .B(n_491), .CI(n_490), .CO(n_85), .S(n_84));
   FA_X1 i_403 (.A(n_59), .B(n_57), .CI(n_489), .CO(n_87), .S(n_86));
   FA_X1 i_404 (.A(n_488), .B(n_487), .CI(n_486), .CO(n_89), .S(n_88));
   FA_X1 i_405 (.A(n_485), .B(n_484), .CI(n_483), .CO(n_91), .S(n_90));
   FA_X1 i_406 (.A(n_61), .B(n_84), .CI(n_82), .CO(n_93), .S(n_92));
   FA_X1 i_407 (.A(n_65), .B(n_63), .CI(n_86), .CO(n_95), .S(n_94));
   FA_X1 i_408 (.A(n_69), .B(n_67), .CI(n_90), .CO(n_97), .S(n_96));
   FA_X1 i_409 (.A(n_88), .B(n_71), .CI(n_94), .CO(n_99), .S(n_98));
   FA_X1 i_410 (.A(n_92), .B(n_73), .CI(n_96), .CO(n_101), .S(n_100));
   FA_X1 i_411 (.A(n_75), .B(n_98), .CI(n_77), .CO(n_103), .S(n_102));
   FA_X1 i_412 (.A(n_100), .B(n_79), .CI(n_102), .CO(n_105), .S(n_104));
   FA_X1 i_413 (.A(n_482), .B(n_481), .CI(n_480), .CO(n_107), .S(n_106));
   FA_X1 i_414 (.A(n_479), .B(n_478), .CI(n_477), .CO(n_109), .S(n_108));
   FA_X1 i_415 (.A(n_476), .B(n_85), .CI(n_83), .CO(n_111), .S(n_110));
   FA_X1 i_416 (.A(n_2084), .B(n_474), .CI(n_473), .CO(n_113), .S(n_112));
   FA_X1 i_417 (.A(n_472), .B(n_471), .CI(n_470), .CO(n_115), .S(n_114));
   FA_X1 i_418 (.A(n_469), .B(n_108), .CI(n_106), .CO(n_117), .S(n_116));
   FA_X1 i_419 (.A(n_91), .B(n_89), .CI(n_87), .CO(n_119), .S(n_118));
   FA_X1 i_420 (.A(n_110), .B(n_93), .CI(n_114), .CO(n_121), .S(n_120));
   FA_X1 i_421 (.A(n_112), .B(n_95), .CI(n_118), .CO(n_123), .S(n_122));
   FA_X1 i_422 (.A(n_116), .B(n_97), .CI(n_120), .CO(n_125), .S(n_124));
   FA_X1 i_423 (.A(n_99), .B(n_122), .CI(n_101), .CO(n_127), .S(n_126));
   FA_X1 i_424 (.A(n_124), .B(n_103), .CI(n_126), .CO(n_129), .S(n_128));
   FA_X1 i_425 (.A(n_468), .B(n_467), .CI(n_466), .CO(n_131), .S(n_130));
   FA_X1 i_426 (.A(n_465), .B(n_464), .CI(n_463), .CO(n_133), .S(n_132));
   FA_X1 i_427 (.A(n_109), .B(n_107), .CI(n_462), .CO(n_135), .S(n_134));
   FA_X1 i_428 (.A(n_461), .B(n_460), .CI(n_459), .CO(n_137), .S(n_136));
   FA_X1 i_429 (.A(n_458), .B(n_457), .CI(n_111), .CO(n_139), .S(n_138));
   FA_X1 i_430 (.A(n_132), .B(n_130), .CI(n_115), .CO(n_141), .S(n_140));
   FA_X1 i_431 (.A(n_113), .B(n_134), .CI(n_119), .CO(n_143), .S(n_142));
   FA_X1 i_432 (.A(n_117), .B(n_138), .CI(n_136), .CO(n_145), .S(n_144));
   FA_X1 i_433 (.A(n_140), .B(n_121), .CI(n_142), .CO(n_147), .S(n_146));
   FA_X1 i_434 (.A(n_123), .B(n_144), .CI(n_125), .CO(n_149), .S(n_148));
   FA_X1 i_435 (.A(n_146), .B(n_127), .CI(n_148), .CO(n_151), .S(n_150));
   FA_X1 i_436 (.A(n_456), .B(n_455), .CI(n_454), .CO(n_153), .S(n_152));
   FA_X1 i_437 (.A(n_453), .B(n_452), .CI(n_133), .CO(n_155), .S(n_154));
   FA_X1 i_438 (.A(n_131), .B(n_451), .CI(n_450), .CO(n_157), .S(n_156));
   FA_X1 i_439 (.A(n_449), .B(n_448), .CI(n_447), .CO(n_159), .S(n_158));
   FA_X1 i_440 (.A(n_446), .B(n_154), .CI(n_152), .CO(n_161), .S(n_160));
   FA_X1 i_441 (.A(n_137), .B(n_135), .CI(n_139), .CO(n_163), .S(n_162));
   FA_X1 i_442 (.A(n_141), .B(n_158), .CI(n_156), .CO(n_165), .S(n_164));
   FA_X1 i_443 (.A(n_143), .B(n_162), .CI(n_160), .CO(n_167), .S(n_166));
   FA_X1 i_444 (.A(n_145), .B(n_164), .CI(n_147), .CO(n_169), .S(n_168));
   FA_X1 i_445 (.A(n_166), .B(n_149), .CI(n_168), .CO(n_171), .S(n_170));
   FA_X1 i_446 (.A(n_543), .B(n_445), .CI(n_444), .CO(n_173), .S(n_172));
   FA_X1 i_447 (.A(n_443), .B(n_442), .CI(n_441), .CO(n_175), .S(n_174));
   FA_X1 i_448 (.A(n_153), .B(n_440), .CI(n_439), .CO(n_177), .S(n_176));
   FA_X1 i_449 (.A(n_438), .B(n_437), .CI(n_436), .CO(n_179), .S(n_178));
   FA_X1 i_450 (.A(n_435), .B(n_155), .CI(n_174), .CO(n_181), .S(n_180));
   FA_X1 i_451 (.A(n_172), .B(n_159), .CI(n_157), .CO(n_183), .S(n_182));
   FA_X1 i_452 (.A(n_176), .B(n_161), .CI(n_163), .CO(n_185), .S(n_184));
   FA_X1 i_453 (.A(n_178), .B(n_180), .CI(n_182), .CO(n_187), .S(n_186));
   FA_X1 i_454 (.A(n_165), .B(n_184), .CI(n_167), .CO(n_189), .S(n_188));
   FA_X1 i_455 (.A(n_186), .B(n_169), .CI(n_188), .CO(n_191), .S(n_190));
   FA_X1 i_456 (.A(n_434), .B(n_433), .CI(n_432), .CO(n_193), .S(n_192));
   FA_X1 i_457 (.A(n_431), .B(n_430), .CI(n_175), .CO(n_195), .S(n_194));
   FA_X1 i_458 (.A(n_173), .B(n_429), .CI(n_428), .CO(n_197), .S(n_196));
   FA_X1 i_459 (.A(n_427), .B(n_426), .CI(n_425), .CO(n_199), .S(n_198));
   FA_X1 i_460 (.A(n_194), .B(n_192), .CI(n_179), .CO(n_201), .S(n_200));
   FA_X1 i_461 (.A(n_177), .B(n_183), .CI(n_181), .CO(n_203), .S(n_202));
   FA_X1 i_462 (.A(n_198), .B(n_196), .CI(n_185), .CO(n_205), .S(n_204));
   FA_X1 i_463 (.A(n_200), .B(n_202), .CI(n_187), .CO(n_207), .S(n_206));
   FA_X1 i_464 (.A(n_204), .B(n_189), .CI(n_206), .CO(n_209), .S(n_208));
   FA_X1 i_465 (.A(n_424), .B(n_423), .CI(n_422), .CO(n_211), .S(n_210));
   FA_X1 i_466 (.A(n_421), .B(n_193), .CI(n_420), .CO(n_213), .S(n_212));
   FA_X1 i_467 (.A(n_419), .B(n_418), .CI(n_417), .CO(n_215), .S(n_214));
   FA_X1 i_468 (.A(n_416), .B(n_195), .CI(n_210), .CO(n_217), .S(n_216));
   FA_X1 i_469 (.A(n_199), .B(n_197), .CI(n_212), .CO(n_219), .S(n_218));
   FA_X1 i_470 (.A(n_201), .B(n_214), .CI(n_216), .CO(n_221), .S(n_220));
   FA_X1 i_471 (.A(n_203), .B(n_218), .CI(n_205), .CO(n_223), .S(n_222));
   FA_X1 i_472 (.A(n_220), .B(n_207), .CI(n_222), .CO(n_225), .S(n_224));
   FA_X1 i_473 (.A(n_639), .B(n_415), .CI(n_414), .CO(n_227), .S(n_226));
   FA_X1 i_474 (.A(n_413), .B(n_412), .CI(n_211), .CO(n_229), .S(n_228));
   FA_X1 i_475 (.A(n_2263), .B(n_410), .CI(n_409), .CO(n_231), .S(n_230));
   FA_X1 i_476 (.A(n_408), .B(n_407), .CI(n_228), .CO(n_233), .S(n_232));
   FA_X1 i_477 (.A(n_226), .B(n_215), .CI(n_213), .CO(n_235), .S(n_234));
   FA_X1 i_478 (.A(n_217), .B(n_232), .CI(n_230), .CO(n_237), .S(n_236));
   FA_X1 i_479 (.A(n_219), .B(n_234), .CI(n_221), .CO(n_239), .S(n_238));
   FA_X1 i_480 (.A(n_223), .B(n_236), .CI(n_238), .CO(n_241), .S(n_240));
   FA_X1 i_481 (.A(n_403), .B(n_227), .CI(n_402), .CO(n_243), .S(n_242));
   FA_X1 i_482 (.A(n_401), .B(n_400), .CI(n_399), .CO(n_245), .S(n_244));
   FA_X1 i_483 (.A(n_229), .B(n_2865), .CI(n_231), .CO(n_247), .S(n_246));
   FA_X1 i_484 (.A(n_242), .B(n_235), .CI(n_233), .CO(n_249), .S(n_248));
   FA_X1 i_485 (.A(n_244), .B(n_246), .CI(n_237), .CO(n_251), .S(n_250));
   FA_X1 i_486 (.A(n_248), .B(n_239), .CI(n_250), .CO(n_253), .S(n_252));
   FA_X1 i_487 (.A(n_393), .B(n_392), .CI(n_2966), .CO(n_255), .S(n_254));
   FA_X1 i_488 (.A(n_245), .B(n_243), .CI(n_247), .CO(n_257), .S(n_256));
   FA_X1 i_489 (.A(n_254), .B(n_2893), .CI(n_249), .CO(n_259), .S(n_258));
   FA_X1 i_490 (.A(n_256), .B(n_251), .CI(n_258), .CO(n_261), .S(n_260));
   FA_X1 i_491 (.A(n_390), .B(n_389), .CI(n_388), .CO(n_263), .S(n_262));
   FA_X1 i_492 (.A(n_255), .B(n_262), .CI(n_257), .CO(n_265), .S(n_264));
   FA_X1 i_493 (.A(n_2978), .B(n_259), .CI(n_264), .CO(n_267), .S(n_266));
   FA_X1 i_494 (.A(n_387), .B(n_386), .CI(n_385), .CO(n_269), .S(n_268));
   FA_X1 i_495 (.A(n_2863), .B(n_384), .CI(n_383), .CO(n_271), .S(n_270));
   FA_X1 i_496 (.A(n_382), .B(n_2972), .CI(n_268), .CO(n_273), .S(n_272));
   FA_X1 i_497 (.A(n_263), .B(n_270), .CI(n_272), .CO(n_275), .S(n_274));
   FA_X1 i_498 (.A(n_2980), .B(n_265), .CI(n_274), .CO(n_277), .S(n_276));
   FA_X1 i_499 (.A(n_381), .B(n_380), .CI(n_269), .CO(n_279), .S(n_278));
   FA_X1 i_500 (.A(n_379), .B(n_378), .CI(n_377), .CO(n_281), .S(n_280));
   FA_X1 i_501 (.A(n_278), .B(n_271), .CI(n_273), .CO(n_283), .S(n_282));
   FA_X1 i_502 (.A(n_280), .B(n_282), .CI(n_275), .CO(n_285), .S(n_284));
   FA_X1 i_503 (.A(n_831), .B(n_376), .CI(n_375), .CO(n_287), .S(n_286));
   FA_X1 i_504 (.A(n_3579), .B(n_374), .CI(n_373), .CO(n_289), .S(n_288));
   FA_X1 i_505 (.A(n_279), .B(n_286), .CI(n_281), .CO(n_291), .S(n_290));
   FA_X1 i_506 (.A(n_288), .B(n_283), .CI(n_290), .CO(n_293), .S(n_292));
   FA_X1 i_507 (.A(n_372), .B(n_371), .CI(n_287), .CO(n_295), .S(n_294));
   FA_X1 i_508 (.A(n_370), .B(n_369), .CI(n_294), .CO(n_297), .S(n_296));
   FA_X1 i_509 (.A(n_289), .B(n_291), .CI(n_296), .CO(n_299), .S(n_298));
   FA_X1 i_510 (.A(n_295), .B(n_297), .CI(n_3651), .CO(n_301), .S(n_300));
   FA_X1 i_511 (.A(n_368), .B(n_367), .CI(n_3650), .CO(n_303), .S(n_302));
   FA_X1 i_512 (.A(n_1022), .B(n_991), .CI(n_366), .CO(n_305), .S(n_304));
   FA_X1 i_4122 (.A(n_1034), .B(n_1029), .CI(n_365), .CO(n_306), .S(out[3]));
   FA_X1 i_4123 (.A(n_1039), .B(n_1052), .CI(n_306), .CO(n_307), .S(out[4]));
   FA_X1 i_4124 (.A(n_1070), .B(n_1068), .CI(n_307), .CO(n_308), .S(out[5]));
   FA_X1 i_4125 (.A(n_1096), .B(n_601), .CI(n_308), .CO(n_309), .S(out[6]));
   FA_X1 i_4126 (.A(n_1122), .B(n_602), .CI(n_309), .CO(n_310), .S(out[7]));
   FA_X1 i_4127 (.A(n_1151), .B(n_1153), .CI(n_310), .CO(n_311), .S(out[8]));
   FA_X1 i_4128 (.A(n_1190), .B(n_1188), .CI(n_311), .CO(n_312), .S(out[9]));
   FA_X1 i_4129 (.A(n_1229), .B(n_1227), .CI(n_312), .CO(n_313), .S(out[10]));
   FA_X1 i_4130 (.A(n_1267), .B(n_1269), .CI(n_313), .CO(n_314), .S(out[11]));
   FA_X1 i_4131 (.A(n_1315), .B(n_1317), .CI(n_314), .CO(n_315), .S(out[12]));
   FA_X1 i_513 (.A(n_1365), .B(n_1367), .CI(n_315), .CO(n_316), .S(out[13]));
   FA_X1 i_514 (.A(n_1416), .B(n_1418), .CI(n_316), .CO(n_317), .S(out[14]));
   FA_X1 i_515 (.A(n_1475), .B(n_1477), .CI(n_317), .CO(n_318), .S(out[15]));
   FA_X1 i_516 (.A(n_1536), .B(n_1538), .CI(n_318), .CO(n_319), .S(out[16]));
   FA_X1 i_517 (.A(n_1598), .B(n_1600), .CI(n_319), .CO(n_320), .S(out[17]));
   FA_X1 i_518 (.A(n_1601), .B(n_1670), .CI(n_320), .CO(n_321), .S(out[18]));
   FA_X1 i_519 (.A(n_1671), .B(n_1742), .CI(n_321), .CO(n_322), .S(out[19]));
   FA_X1 i_520 (.A(n_1813), .B(n_1815), .CI(n_322), .CO(n_323), .S(out[20]));
   FA_X1 i_521 (.A(n_1816), .B(n_1896), .CI(n_323), .CO(n_324), .S(out[21]));
   FA_X1 i_522 (.A(n_1897), .B(n_1979), .CI(n_324), .CO(n_325), .S(out[22]));
   FA_X1 i_523 (.A(n_1980), .B(n_2063), .CI(n_325), .CO(n_326), .S(out[23]));
   FA_X1 i_524 (.A(n_2064), .B(n_2155), .CI(n_326), .CO(n_327), .S(out[24]));
   FA_X1 i_525 (.A(n_2247), .B(n_2249), .CI(n_327), .CO(n_328), .S(out[25]));
   FA_X1 i_526 (.A(n_2250), .B(n_2344), .CI(n_328), .CO(n_329), .S(out[26]));
   FA_X1 i_527 (.A(n_2345), .B(n_2447), .CI(n_329), .CO(n_330), .S(out[27]));
   FA_X1 i_528 (.A(n_2448), .B(n_2552), .CI(n_330), .CO(n_331), .S(out[28]));
   FA_X1 i_529 (.A(n_2553), .B(n_2658), .CI(n_331), .CO(n_332), .S(out[29]));
   FA_X1 i_530 (.A(n_2659), .B(n_2772), .CI(n_332), .CO(n_333), .S(out[30]));
   FA_X1 i_531 (.A(n_2773), .B(n_2889), .CI(n_333), .CO(n_334), .S(out[31]));
   FA_X1 i_532 (.A(n_2890), .B(n_3002), .CI(n_334), .CO(n_335), .S(out[32]));
   FA_X1 i_533 (.A(n_3003), .B(n_3112), .CI(n_335), .CO(n_336), .S(out[33]));
   FA_X1 i_534 (.A(n_3113), .B(n_3220), .CI(n_336), .CO(n_337), .S(out[34]));
   FA_X1 i_535 (.A(n_3320), .B(n_3221), .CI(n_337), .CO(n_338), .S(out[35]));
   FA_X1 i_536 (.A(n_3321), .B(n_3419), .CI(n_338), .CO(n_339), .S(out[36]));
   FA_X1 i_537 (.A(n_3420), .B(n_3516), .CI(n_339), .CO(n_340), .S(out[37]));
   FA_X1 i_538 (.A(n_3517), .B(n_3605), .CI(n_340), .CO(n_341), .S(out[38]));
   FA_X1 i_539 (.A(n_3606), .B(n_3693), .CI(n_341), .CO(n_342), .S(out[39]));
   FA_X1 i_540 (.A(n_3694), .B(n_26), .CI(n_342), .CO(n_343), .S(out[40]));
   FA_X1 i_541 (.A(n_27), .B(n_54), .CI(n_343), .CO(n_344), .S(out[41]));
   FA_X1 i_542 (.A(n_55), .B(n_80), .CI(n_344), .CO(n_345), .S(out[42]));
   FA_X1 i_543 (.A(n_81), .B(n_104), .CI(n_345), .CO(n_346), .S(out[43]));
   FA_X1 i_544 (.A(n_105), .B(n_128), .CI(n_346), .CO(n_347), .S(out[44]));
   FA_X1 i_545 (.A(n_129), .B(n_150), .CI(n_347), .CO(n_348), .S(out[45]));
   FA_X1 i_546 (.A(n_151), .B(n_170), .CI(n_348), .CO(n_349), .S(out[46]));
   FA_X1 i_547 (.A(n_171), .B(n_190), .CI(n_349), .CO(n_350), .S(out[47]));
   FA_X1 i_548 (.A(n_191), .B(n_208), .CI(n_350), .CO(n_351), .S(out[48]));
   FA_X1 i_549 (.A(n_224), .B(n_209), .CI(n_351), .CO(n_352), .S(out[49]));
   FA_X1 i_550 (.A(n_225), .B(n_240), .CI(n_352), .CO(n_353), .S(out[50]));
   FA_X1 i_551 (.A(n_241), .B(n_252), .CI(n_353), .CO(n_354), .S(out[51]));
   FA_X1 i_552 (.A(n_260), .B(n_253), .CI(n_354), .CO(n_355), .S(out[52]));
   FA_X1 i_553 (.A(n_261), .B(n_266), .CI(n_355), .CO(n_356), .S(out[53]));
   FA_X1 i_554 (.A(n_267), .B(n_276), .CI(n_356), .CO(n_357), .S(out[54]));
   FA_X1 i_555 (.A(n_284), .B(n_277), .CI(n_357), .CO(n_358), .S(out[55]));
   FA_X1 i_556 (.A(n_285), .B(n_292), .CI(n_358), .CO(n_359), .S(out[56]));
   FA_X1 i_557 (.A(n_298), .B(n_293), .CI(n_359), .CO(n_360), .S(out[57]));
   FA_X1 i_558 (.A(n_299), .B(n_300), .CI(n_360), .CO(n_361), .S(out[58]));
   FA_X1 i_559 (.A(n_3654), .B(n_301), .CI(n_361), .CO(n_362), .S(out[59]));
   FA_X1 i_560 (.A(n_3655), .B(n_302), .CI(n_362), .CO(n_363), .S(out[60]));
   FA_X1 i_561 (.A(n_304), .B(n_303), .CI(n_363), .CO(n_364), .S(out[61]));
   NAND2_X1 i_562 (.A1(in2[2]), .A2(in1[1]), .ZN(n_518));
   NOR2_X1 i_563 (.A1(n_518), .A2(n_679), .ZN(n_520));
   AOI22_X1 i_564 (.A1(in2[2]), .A2(in1[2]), .B1(in2[3]), .B2(in1[1]), .ZN(n_521));
   NOR2_X1 i_4 (.A1(n_520), .A2(n_521), .ZN(n_522));
   NAND2_X1 i_565 (.A1(in2[4]), .A2(in1[0]), .ZN(n_523));
   XNOR2_X1 i_6 (.A(n_522), .B(n_523), .ZN(n_1039));
   NOR2_X1 i_566 (.A1(n_690), .A2(n_692), .ZN(out[0]));
   NOR3_X1 i_567 (.A1(n_518), .A2(n_1377), .A3(n_690), .ZN(n_527));
   AOI22_X1 i_568 (.A1(in2[1]), .A2(in1[1]), .B1(in2[2]), .B2(in1[0]), .ZN(n_528));
   NOR2_X1 i_569 (.A1(n_527), .A2(n_528), .ZN(n_529));
   AOI21_X1 i_570 (.A(n_529), .B1(in1[2]), .B2(in2[0]), .ZN(n_530));
   NAND3_X1 i_571 (.A1(out[0]), .A2(in2[1]), .A3(in1[1]), .ZN(n_531));
   NAND3_X1 i_572 (.A1(n_529), .A2(in1[2]), .A3(in2[0]), .ZN(n_532));
   AOI21_X1 i_17 (.A(n_530), .B1(n_531), .B2(n_532), .ZN(n_365));
   INV_X1 i_573 (.A(n_518), .ZN(n_533));
   NAND3_X1 i_574 (.A1(n_533), .A2(in1[2]), .A3(in2[1]), .ZN(n_534));
   AOI21_X1 i_575 (.A(n_533), .B1(in1[2]), .B2(in2[1]), .ZN(n_535));
   INV_X1 i_21 (.A(n_535), .ZN(n_536));
   NAND2_X1 i_22 (.A1(n_534), .A2(n_536), .ZN(n_537));
   NAND2_X1 i_576 (.A1(in2[3]), .A2(in1[0]), .ZN(n_538));
   XOR2_X1 i_24 (.A(n_537), .B(n_538), .Z(n_1029));
   AND2_X1 i_577 (.A1(in1[3]), .A2(in2[0]), .ZN(n_539));
   XOR2_X1 i_26 (.A(n_527), .B(n_539), .Z(n_1034));
   NOR2_X1 i_578 (.A1(n_1382), .A2(n_1602), .ZN(n_542));
   XOR2_X1 i_579 (.A(n_542), .B(n_3730), .Z(n_545));
   NOR2_X1 i_580 (.A1(n_1384), .A2(n_1581), .ZN(n_548));
   AOI22_X1 i_581 (.A1(n_545), .A2(n_548), .B1(n_542), .B2(n_3730), .ZN(n_366));
   NAND2_X1 i_582 (.A1(in1[31]), .A2(in2[30]), .ZN(n_991));
   NAND2_X1 i_583 (.A1(in2[31]), .A2(in1[30]), .ZN(n_1022));
   XNOR2_X1 i_584 (.A(n_545), .B(n_548), .ZN(n_367));
   INV_X1 i_585 (.A(n_3728), .ZN(n_552));
   AOI21_X1 i_586 (.A(n_3725), .B1(n_552), .B2(n_3724), .ZN(n_368));
   INV_X1 i_587 (.A(n_3715), .ZN(n_580));
   NAND2_X1 i_588 (.A1(n_3716), .A2(n_580), .ZN(n_581));
   XOR2_X1 i_589 (.A(n_581), .B(n_3714), .Z(n_369));
   NAND2_X1 i_590 (.A1(n_3723), .A2(n_3722), .ZN(n_582));
   XOR2_X1 i_591 (.A(n_582), .B(n_3718), .Z(n_370));
   NAND3_X1 i_592 (.A1(n_3717), .A2(in2[29]), .A3(in1[26]), .ZN(n_583));
   AOI22_X1 i_593 (.A1(in2[30]), .A2(in1[26]), .B1(in2[29]), .B2(in1[27]), 
      .ZN(n_584));
   AND2_X1 i_594 (.A1(in2[31]), .A2(in1[25]), .ZN(n_585));
   OAI21_X1 i_595 (.A(n_583), .B1(n_584), .B2(n_585), .ZN(n_371));
   NAND4_X1 i_596 (.A1(in1[29]), .A2(in1[30]), .A3(in2[27]), .A4(in2[26]), 
      .ZN(n_586));
   AOI22_X1 i_597 (.A1(in1[29]), .A2(in2[27]), .B1(in1[30]), .B2(in2[26]), 
      .ZN(n_587));
   NAND2_X1 i_598 (.A1(in1[28]), .A2(in2[28]), .ZN(n_588));
   OAI21_X1 i_599 (.A(n_586), .B1(n_587), .B2(n_588), .ZN(n_372));
   INV_X1 i_600 (.A(n_584), .ZN(n_589));
   NAND2_X1 i_601 (.A1(n_583), .A2(n_589), .ZN(n_590));
   XOR2_X1 i_602 (.A(n_590), .B(n_585), .Z(n_373));
   INV_X1 i_603 (.A(n_587), .ZN(n_591));
   NAND2_X1 i_604 (.A1(n_591), .A2(n_586), .ZN(n_592));
   XOR2_X1 i_605 (.A(n_592), .B(n_588), .Z(n_374));
   NAND4_X1 i_606 (.A1(in2[30]), .A2(in2[29]), .A3(in1[26]), .A4(in1[25]), 
      .ZN(n_605));
   AOI22_X1 i_607 (.A1(in2[30]), .A2(in1[25]), .B1(in2[29]), .B2(in1[26]), 
      .ZN(n_606));
   AND2_X1 i_608 (.A1(in2[31]), .A2(in1[24]), .ZN(n_607));
   OAI21_X1 i_609 (.A(n_605), .B1(n_606), .B2(n_607), .ZN(n_375));
   NOR2_X1 i_610 (.A1(n_1580), .A2(n_3732), .ZN(n_608));
   NAND3_X1 i_611 (.A1(n_608), .A2(in1[29]), .A3(in2[26]), .ZN(n_609));
   AOI21_X1 i_612 (.A(n_608), .B1(in1[29]), .B2(in2[26]), .ZN(n_610));
   NAND2_X1 i_613 (.A1(in2[28]), .A2(in1[27]), .ZN(n_611));
   OAI21_X1 i_614 (.A(n_609), .B1(n_610), .B2(n_611), .ZN(n_376));
   NAND2_X1 i_615 (.A1(in1[31]), .A2(in2[25]), .ZN(n_831));
   INV_X1 i_616 (.A(n_606), .ZN(n_612));
   NAND2_X1 i_617 (.A1(n_612), .A2(n_605), .ZN(n_613));
   XOR2_X1 i_618 (.A(n_613), .B(n_607), .Z(n_377));
   INV_X1 i_619 (.A(n_610), .ZN(n_614));
   NAND2_X1 i_620 (.A1(n_609), .A2(n_614), .ZN(n_615));
   XOR2_X1 i_621 (.A(n_615), .B(n_611), .Z(n_378));
   XNOR2_X1 i_622 (.A(n_3607), .B(n_3621), .ZN(n_379));
   NAND4_X1 i_623 (.A1(in2[30]), .A2(in2[29]), .A3(in1[25]), .A4(in1[24]), 
      .ZN(n_616));
   AOI22_X1 i_624 (.A1(in2[30]), .A2(in1[24]), .B1(in2[29]), .B2(in1[25]), 
      .ZN(n_617));
   AND2_X1 i_625 (.A1(in2[31]), .A2(in1[23]), .ZN(n_618));
   OAI21_X1 i_626 (.A(n_616), .B1(n_617), .B2(n_618), .ZN(n_380));
   NAND4_X1 i_627 (.A1(in1[28]), .A2(in1[27]), .A3(in2[27]), .A4(in2[26]), 
      .ZN(n_619));
   AOI22_X1 i_628 (.A1(in1[27]), .A2(in2[27]), .B1(in1[28]), .B2(in2[26]), 
      .ZN(n_620));
   NAND2_X1 i_629 (.A1(in2[28]), .A2(in1[26]), .ZN(n_621));
   OAI21_X1 i_630 (.A(n_619), .B1(n_620), .B2(n_621), .ZN(n_381));
   INV_X1 i_631 (.A(n_617), .ZN(n_622));
   NAND2_X1 i_632 (.A1(n_622), .A2(n_616), .ZN(n_623));
   XOR2_X1 i_633 (.A(n_623), .B(n_618), .Z(n_382));
   INV_X1 i_634 (.A(n_620), .ZN(n_624));
   NAND2_X1 i_635 (.A1(n_624), .A2(n_619), .ZN(n_625));
   XOR2_X1 i_636 (.A(n_625), .B(n_621), .Z(n_383));
   NAND2_X1 i_637 (.A1(n_3648), .A2(n_3647), .ZN(n_626));
   XOR2_X1 i_638 (.A(n_626), .B(n_3643), .Z(n_384));
   NAND4_X1 i_639 (.A1(in2[30]), .A2(in2[29]), .A3(in1[23]), .A4(in1[24]), 
      .ZN(n_627));
   AOI22_X1 i_640 (.A1(in2[30]), .A2(in1[23]), .B1(in2[29]), .B2(in1[24]), 
      .ZN(n_628));
   AND2_X1 i_641 (.A1(in2[31]), .A2(in1[22]), .ZN(n_629));
   OAI21_X1 i_642 (.A(n_627), .B1(n_628), .B2(n_629), .ZN(n_385));
   NAND4_X1 i_643 (.A1(in1[26]), .A2(in1[27]), .A3(in2[27]), .A4(in2[26]), 
      .ZN(n_630));
   AOI22_X1 i_644 (.A1(in1[26]), .A2(in2[27]), .B1(in1[27]), .B2(in2[26]), 
      .ZN(n_631));
   NAND2_X1 i_645 (.A1(in2[28]), .A2(in1[25]), .ZN(n_632));
   OAI21_X1 i_646 (.A(n_630), .B1(n_631), .B2(n_632), .ZN(n_386));
   NAND4_X1 i_647 (.A1(in1[29]), .A2(in1[30]), .A3(in2[24]), .A4(in2[23]), 
      .ZN(n_633));
   AOI22_X1 i_648 (.A1(in1[29]), .A2(in2[24]), .B1(in1[30]), .B2(in2[23]), 
      .ZN(n_634));
   NAND2_X1 i_649 (.A1(in1[28]), .A2(in2[25]), .ZN(n_635));
   OAI21_X1 i_650 (.A(n_633), .B1(n_634), .B2(n_635), .ZN(n_387));
   INV_X1 i_651 (.A(n_628), .ZN(n_636));
   NAND2_X1 i_652 (.A1(n_636), .A2(n_627), .ZN(n_637));
   XOR2_X1 i_653 (.A(n_637), .B(n_629), .Z(n_388));
   INV_X1 i_654 (.A(n_631), .ZN(n_638));
   NAND2_X1 i_655 (.A1(n_638), .A2(n_630), .ZN(n_640));
   XOR2_X1 i_656 (.A(n_640), .B(n_632), .Z(n_389));
   INV_X1 i_657 (.A(n_634), .ZN(n_641));
   NAND2_X1 i_658 (.A1(n_641), .A2(n_633), .ZN(n_642));
   XOR2_X1 i_659 (.A(n_642), .B(n_635), .Z(n_390));
   INV_X1 i_660 (.A(n_3291), .ZN(n_665));
   NAND2_X1 i_661 (.A1(n_665), .A2(n_3292), .ZN(n_666));
   XOR2_X1 i_662 (.A(n_666), .B(n_3289), .Z(n_392));
   INV_X1 i_663 (.A(n_3568), .ZN(n_667));
   NAND2_X1 i_664 (.A1(n_667), .A2(n_3569), .ZN(n_668));
   XOR2_X1 i_665 (.A(n_668), .B(n_3567), .Z(n_393));
   INV_X1 i_666 (.A(n_3203), .ZN(n_680));
   NAND2_X1 i_667 (.A1(n_680), .A2(n_3205), .ZN(n_681));
   XOR2_X1 i_668 (.A(n_681), .B(n_3193), .Z(n_399));
   INV_X1 i_669 (.A(n_3207), .ZN(n_682));
   NAND2_X1 i_670 (.A1(n_682), .A2(n_3208), .ZN(n_683));
   XOR2_X1 i_671 (.A(n_683), .B(n_3206), .Z(n_400));
   INV_X1 i_672 (.A(n_3213), .ZN(n_684));
   NAND2_X1 i_673 (.A1(n_684), .A2(n_3287), .ZN(n_685));
   XOR2_X1 i_674 (.A(n_685), .B(n_3212), .Z(n_401));
   NAND2_X1 i_675 (.A1(n_3313), .A2(n_3312), .ZN(n_686));
   XOR2_X1 i_676 (.A(n_686), .B(n_3303), .Z(n_402));
   NAND4_X1 i_677 (.A1(in2[30]), .A2(in2[29]), .A3(in1[20]), .A4(in1[21]), 
      .ZN(n_687));
   AOI22_X1 i_678 (.A1(in2[30]), .A2(in1[20]), .B1(in2[29]), .B2(in1[21]), 
      .ZN(n_688));
   AND2_X1 i_679 (.A1(in2[31]), .A2(in1[19]), .ZN(n_689));
   OAI21_X1 i_680 (.A(n_687), .B1(n_688), .B2(n_689), .ZN(n_403));
   INV_X1 i_681 (.A(n_688), .ZN(n_699));
   NAND2_X1 i_682 (.A1(n_699), .A2(n_687), .ZN(n_700));
   XOR2_X1 i_683 (.A(n_700), .B(n_689), .Z(n_407));
   INV_X1 i_684 (.A(n_3392), .ZN(n_701));
   NAND2_X1 i_685 (.A1(n_701), .A2(n_3401), .ZN(n_702));
   XOR2_X1 i_686 (.A(n_702), .B(n_3390), .Z(n_408));
   INV_X1 i_687 (.A(n_3486), .ZN(n_703));
   NAND2_X1 i_688 (.A1(n_703), .A2(n_3488), .ZN(n_704));
   XOR2_X1 i_689 (.A(n_704), .B(n_3402), .Z(n_409));
   INV_X1 i_690 (.A(n_3565), .ZN(n_705));
   NAND2_X1 i_691 (.A1(n_705), .A2(n_3566), .ZN(n_706));
   XOR2_X1 i_692 (.A(n_706), .B(n_3562), .Z(n_410));
   NAND4_X1 i_693 (.A1(in2[30]), .A2(in2[29]), .A3(in1[20]), .A4(in1[19]), 
      .ZN(n_719));
   AOI22_X1 i_694 (.A1(in2[30]), .A2(in1[19]), .B1(in2[29]), .B2(in1[20]), 
      .ZN(n_720));
   AND2_X1 i_695 (.A1(in2[31]), .A2(in1[18]), .ZN(n_721));
   OAI21_X1 i_696 (.A(n_719), .B1(n_720), .B2(n_721), .ZN(n_412));
   NAND4_X1 i_697 (.A1(in2[27]), .A2(in2[26]), .A3(in1[23]), .A4(in1[22]), 
      .ZN(n_722));
   AOI22_X1 i_698 (.A1(in2[27]), .A2(in1[22]), .B1(in2[26]), .B2(in1[23]), 
      .ZN(n_723));
   NAND2_X1 i_699 (.A1(in2[28]), .A2(in1[21]), .ZN(n_724));
   OAI21_X1 i_700 (.A(n_722), .B1(n_723), .B2(n_724), .ZN(n_413));
   NAND4_X1 i_701 (.A1(in1[26]), .A2(in1[25]), .A3(in2[24]), .A4(in2[23]), 
      .ZN(n_725));
   AOI22_X1 i_702 (.A1(in1[25]), .A2(in2[24]), .B1(in1[26]), .B2(in2[23]), 
      .ZN(n_726));
   NAND2_X1 i_703 (.A1(in2[25]), .A2(in1[24]), .ZN(n_727));
   OAI21_X1 i_704 (.A(n_725), .B1(n_726), .B2(n_727), .ZN(n_414));
   NOR2_X1 i_705 (.A1(n_1580), .A2(n_3573), .ZN(n_728));
   NAND3_X1 i_706 (.A1(n_728), .A2(in1[29]), .A3(in2[20]), .ZN(n_729));
   AOI21_X1 i_707 (.A(n_728), .B1(in1[29]), .B2(in2[20]), .ZN(n_730));
   NAND2_X1 i_708 (.A1(in1[27]), .A2(in2[22]), .ZN(n_731));
   OAI21_X1 i_709 (.A(n_729), .B1(n_730), .B2(n_731), .ZN(n_415));
   NAND2_X1 i_710 (.A1(in1[31]), .A2(in2[19]), .ZN(n_639));
   INV_X1 i_711 (.A(n_720), .ZN(n_732));
   NAND2_X1 i_712 (.A1(n_732), .A2(n_719), .ZN(n_733));
   XOR2_X1 i_713 (.A(n_733), .B(n_721), .Z(n_416));
   INV_X1 i_714 (.A(n_723), .ZN(n_734));
   NAND2_X1 i_715 (.A1(n_734), .A2(n_722), .ZN(n_736));
   XOR2_X1 i_716 (.A(n_736), .B(n_724), .Z(n_417));
   INV_X1 i_717 (.A(n_726), .ZN(n_737));
   NAND2_X1 i_718 (.A1(n_737), .A2(n_725), .ZN(n_738));
   XOR2_X1 i_719 (.A(n_738), .B(n_727), .Z(n_418));
   INV_X1 i_720 (.A(n_730), .ZN(n_739));
   NAND2_X1 i_721 (.A1(n_729), .A2(n_739), .ZN(n_740));
   XOR2_X1 i_722 (.A(n_740), .B(n_731), .Z(n_419));
   XNOR2_X1 i_723 (.A(n_2265), .B(n_2305), .ZN(n_420));
   NAND4_X1 i_724 (.A1(in2[30]), .A2(in2[29]), .A3(in1[19]), .A4(in1[18]), 
      .ZN(n_741));
   AOI22_X1 i_725 (.A1(in2[30]), .A2(in1[18]), .B1(in2[29]), .B2(in1[19]), 
      .ZN(n_742));
   AND2_X1 i_726 (.A1(in2[31]), .A2(in1[17]), .ZN(n_743));
   OAI21_X1 i_727 (.A(n_741), .B1(n_742), .B2(n_743), .ZN(n_421));
   NAND4_X1 i_728 (.A1(in2[27]), .A2(in2[26]), .A3(in1[22]), .A4(in1[21]), 
      .ZN(n_744));
   AOI22_X1 i_729 (.A1(in2[27]), .A2(in1[21]), .B1(in2[26]), .B2(in1[22]), 
      .ZN(n_745));
   NAND2_X1 i_730 (.A1(in2[28]), .A2(in1[20]), .ZN(n_746));
   OAI21_X1 i_731 (.A(n_744), .B1(n_745), .B2(n_746), .ZN(n_422));
   NAND4_X1 i_732 (.A1(in1[25]), .A2(in1[24]), .A3(in2[24]), .A4(in2[23]), 
      .ZN(n_747));
   AOI22_X1 i_733 (.A1(in1[24]), .A2(in2[24]), .B1(in1[25]), .B2(in2[23]), 
      .ZN(n_748));
   NAND2_X1 i_734 (.A1(in2[25]), .A2(in1[23]), .ZN(n_749));
   OAI21_X1 i_735 (.A(n_747), .B1(n_748), .B2(n_749), .ZN(n_423));
   NAND4_X1 i_736 (.A1(in1[28]), .A2(in1[27]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_750));
   AOI22_X1 i_737 (.A1(in1[27]), .A2(in2[21]), .B1(in1[28]), .B2(in2[20]), 
      .ZN(n_751));
   NAND2_X1 i_738 (.A1(in1[26]), .A2(in2[22]), .ZN(n_752));
   OAI21_X1 i_739 (.A(n_750), .B1(n_751), .B2(n_752), .ZN(n_424));
   INV_X1 i_740 (.A(n_742), .ZN(n_753));
   NAND2_X1 i_741 (.A1(n_753), .A2(n_741), .ZN(n_754));
   XOR2_X1 i_742 (.A(n_754), .B(n_743), .Z(n_425));
   INV_X1 i_743 (.A(n_745), .ZN(n_755));
   NAND2_X1 i_744 (.A1(n_755), .A2(n_744), .ZN(n_756));
   XOR2_X1 i_745 (.A(n_756), .B(n_746), .Z(n_426));
   INV_X1 i_746 (.A(n_748), .ZN(n_757));
   NAND2_X1 i_747 (.A1(n_757), .A2(n_747), .ZN(n_758));
   XOR2_X1 i_748 (.A(n_758), .B(n_749), .Z(n_427));
   INV_X1 i_749 (.A(n_751), .ZN(n_759));
   NAND2_X1 i_750 (.A1(n_759), .A2(n_750), .ZN(n_760));
   XOR2_X1 i_751 (.A(n_760), .B(n_752), .Z(n_428));
   NAND2_X1 i_752 (.A1(n_2855), .A2(n_2853), .ZN(n_761));
   XOR2_X1 i_753 (.A(n_761), .B(n_2738), .Z(n_429));
   NAND4_X1 i_754 (.A1(in2[30]), .A2(in2[29]), .A3(in1[17]), .A4(in1[18]), 
      .ZN(n_762));
   AOI22_X1 i_755 (.A1(in2[30]), .A2(in1[17]), .B1(in2[29]), .B2(in1[18]), 
      .ZN(n_763));
   AND2_X1 i_756 (.A1(in2[31]), .A2(in1[16]), .ZN(n_764));
   OAI21_X1 i_757 (.A(n_762), .B1(n_763), .B2(n_764), .ZN(n_430));
   NAND4_X1 i_758 (.A1(in2[27]), .A2(in2[26]), .A3(in1[20]), .A4(in1[21]), 
      .ZN(n_765));
   AOI22_X1 i_759 (.A1(in2[27]), .A2(in1[20]), .B1(in2[26]), .B2(in1[21]), 
      .ZN(n_766));
   NAND2_X1 i_760 (.A1(in2[28]), .A2(in1[19]), .ZN(n_767));
   OAI21_X1 i_761 (.A(n_765), .B1(n_766), .B2(n_767), .ZN(n_431));
   NAND4_X1 i_762 (.A1(in1[23]), .A2(in1[24]), .A3(in2[24]), .A4(in2[23]), 
      .ZN(n_768));
   AOI22_X1 i_763 (.A1(in1[23]), .A2(in2[24]), .B1(in1[24]), .B2(in2[23]), 
      .ZN(n_769));
   NAND2_X1 i_764 (.A1(in2[25]), .A2(in1[22]), .ZN(n_770));
   OAI21_X1 i_765 (.A(n_768), .B1(n_769), .B2(n_770), .ZN(n_432));
   NAND4_X1 i_766 (.A1(in1[26]), .A2(in1[27]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_771));
   AOI22_X1 i_767 (.A1(in1[26]), .A2(in2[21]), .B1(in1[27]), .B2(in2[20]), 
      .ZN(n_772));
   NAND2_X1 i_768 (.A1(in1[25]), .A2(in2[22]), .ZN(n_773));
   OAI21_X1 i_769 (.A(n_771), .B1(n_772), .B2(n_773), .ZN(n_433));
   NAND4_X1 i_770 (.A1(in1[29]), .A2(in1[30]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_774));
   AOI22_X1 i_771 (.A1(in1[29]), .A2(in2[18]), .B1(in1[30]), .B2(in2[17]), 
      .ZN(n_775));
   NAND2_X1 i_772 (.A1(in1[28]), .A2(in2[19]), .ZN(n_776));
   OAI21_X1 i_773 (.A(n_774), .B1(n_775), .B2(n_776), .ZN(n_434));
   INV_X1 i_774 (.A(n_763), .ZN(n_777));
   NAND2_X1 i_775 (.A1(n_777), .A2(n_762), .ZN(n_778));
   XOR2_X1 i_776 (.A(n_778), .B(n_764), .Z(n_435));
   INV_X1 i_777 (.A(n_766), .ZN(n_779));
   NAND2_X1 i_778 (.A1(n_779), .A2(n_765), .ZN(n_780));
   XOR2_X1 i_779 (.A(n_780), .B(n_767), .Z(n_436));
   INV_X1 i_780 (.A(n_769), .ZN(n_781));
   NAND2_X1 i_781 (.A1(n_781), .A2(n_768), .ZN(n_782));
   XOR2_X1 i_782 (.A(n_782), .B(n_770), .Z(n_437));
   INV_X1 i_783 (.A(n_772), .ZN(n_783));
   NAND2_X1 i_784 (.A1(n_783), .A2(n_771), .ZN(n_784));
   XOR2_X1 i_785 (.A(n_784), .B(n_773), .Z(n_438));
   INV_X1 i_786 (.A(n_775), .ZN(n_785));
   NAND2_X1 i_787 (.A1(n_785), .A2(n_774), .ZN(n_786));
   XOR2_X1 i_788 (.A(n_786), .B(n_776), .Z(n_439));
   AND2_X1 i_789 (.A1(in1[30]), .A2(in2[16]), .ZN(n_787));
   INV_X1 i_790 (.A(in2[14]), .ZN(n_788));
   OAI211_X1 i_791 (.A(in1[30]), .B(in2[15]), .C1(n_1384), .C2(n_788), .ZN(n_789));
   INV_X1 i_792 (.A(in2[15]), .ZN(n_790));
   OAI211_X1 i_793 (.A(in1[31]), .B(in2[14]), .C1(n_1383), .C2(n_790), .ZN(n_791));
   INV_X1 i_794 (.A(n_791), .ZN(n_792));
   NAND2_X1 i_795 (.A1(in1[29]), .A2(in2[16]), .ZN(n_793));
   OAI21_X1 i_796 (.A(n_789), .B1(n_792), .B2(n_793), .ZN(n_794));
   NOR2_X1 i_797 (.A1(n_1384), .A2(n_790), .ZN(n_795));
   XOR2_X1 i_798 (.A(n_787), .B(n_795), .Z(n_796));
   OAI21_X1 i_799 (.A(n_787), .B1(n_794), .B2(n_796), .ZN(n_797));
   INV_X1 i_800 (.A(n_794), .ZN(n_798));
   OAI21_X1 i_801 (.A(n_797), .B1(n_798), .B2(n_795), .ZN(n_440));
   NAND4_X1 i_802 (.A1(in2[30]), .A2(in2[29]), .A3(in1[17]), .A4(in1[16]), 
      .ZN(n_799));
   AOI22_X1 i_803 (.A1(in2[30]), .A2(in1[16]), .B1(in2[29]), .B2(in1[17]), 
      .ZN(n_800));
   AND2_X1 i_804 (.A1(in2[31]), .A2(in1[15]), .ZN(n_801));
   OAI21_X1 i_805 (.A(n_799), .B1(n_800), .B2(n_801), .ZN(n_441));
   NAND4_X1 i_806 (.A1(in2[27]), .A2(in2[26]), .A3(in1[20]), .A4(in1[19]), 
      .ZN(n_802));
   AOI22_X1 i_807 (.A1(in2[27]), .A2(in1[19]), .B1(in2[26]), .B2(in1[20]), 
      .ZN(n_803));
   NAND2_X1 i_808 (.A1(in2[28]), .A2(in1[18]), .ZN(n_804));
   OAI21_X1 i_809 (.A(n_802), .B1(n_803), .B2(n_804), .ZN(n_442));
   NAND4_X1 i_810 (.A1(in1[23]), .A2(in2[24]), .A3(in2[23]), .A4(in1[22]), 
      .ZN(n_805));
   AOI22_X1 i_811 (.A1(in2[24]), .A2(in1[22]), .B1(in1[23]), .B2(in2[23]), 
      .ZN(n_806));
   NAND2_X1 i_812 (.A1(in2[25]), .A2(in1[21]), .ZN(n_807));
   OAI21_X1 i_813 (.A(n_805), .B1(n_806), .B2(n_807), .ZN(n_443));
   NAND4_X1 i_814 (.A1(in1[26]), .A2(in1[25]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_808));
   AOI22_X1 i_815 (.A1(in1[25]), .A2(in2[21]), .B1(in1[26]), .B2(in2[20]), 
      .ZN(n_809));
   NAND2_X1 i_816 (.A1(in1[24]), .A2(in2[22]), .ZN(n_810));
   OAI21_X1 i_817 (.A(n_808), .B1(n_809), .B2(n_810), .ZN(n_444));
   NOR2_X1 i_818 (.A1(n_1580), .A2(n_2859), .ZN(n_811));
   NAND3_X1 i_819 (.A1(n_811), .A2(in1[29]), .A3(in2[17]), .ZN(n_812));
   AOI21_X1 i_820 (.A(n_811), .B1(in1[29]), .B2(in2[17]), .ZN(n_813));
   NAND2_X1 i_821 (.A1(in1[27]), .A2(in2[19]), .ZN(n_814));
   OAI21_X1 i_822 (.A(n_812), .B1(n_813), .B2(n_814), .ZN(n_445));
   NAND2_X1 i_823 (.A1(in1[31]), .A2(in2[16]), .ZN(n_543));
   INV_X1 i_824 (.A(n_800), .ZN(n_815));
   NAND2_X1 i_825 (.A1(n_815), .A2(n_799), .ZN(n_816));
   XOR2_X1 i_826 (.A(n_816), .B(n_801), .Z(n_446));
   INV_X1 i_827 (.A(n_803), .ZN(n_817));
   NAND2_X1 i_828 (.A1(n_817), .A2(n_802), .ZN(n_818));
   XOR2_X1 i_829 (.A(n_818), .B(n_804), .Z(n_447));
   INV_X1 i_830 (.A(n_806), .ZN(n_819));
   NAND2_X1 i_831 (.A1(n_819), .A2(n_805), .ZN(n_820));
   XOR2_X1 i_832 (.A(n_820), .B(n_807), .Z(n_448));
   INV_X1 i_833 (.A(n_809), .ZN(n_821));
   NAND2_X1 i_834 (.A1(n_821), .A2(n_808), .ZN(n_822));
   XOR2_X1 i_835 (.A(n_822), .B(n_810), .Z(n_449));
   INV_X1 i_836 (.A(n_813), .ZN(n_823));
   NAND2_X1 i_837 (.A1(n_812), .A2(n_823), .ZN(n_824));
   XOR2_X1 i_838 (.A(n_824), .B(n_814), .Z(n_450));
   XNOR2_X1 i_839 (.A(n_796), .B(n_794), .ZN(n_451));
   NAND4_X1 i_840 (.A1(in2[30]), .A2(in2[29]), .A3(in1[16]), .A4(in1[15]), 
      .ZN(n_825));
   AOI22_X1 i_841 (.A1(in2[30]), .A2(in1[15]), .B1(in2[29]), .B2(in1[16]), 
      .ZN(n_826));
   AND2_X1 i_842 (.A1(in2[31]), .A2(in1[14]), .ZN(n_827));
   OAI21_X1 i_843 (.A(n_825), .B1(n_826), .B2(n_827), .ZN(n_452));
   NAND4_X1 i_844 (.A1(in2[27]), .A2(in2[26]), .A3(in1[19]), .A4(in1[18]), 
      .ZN(n_828));
   AOI22_X1 i_845 (.A1(in2[27]), .A2(in1[18]), .B1(in2[26]), .B2(in1[19]), 
      .ZN(n_829));
   NAND2_X1 i_846 (.A1(in2[28]), .A2(in1[17]), .ZN(n_830));
   OAI21_X1 i_847 (.A(n_828), .B1(n_829), .B2(n_830), .ZN(n_453));
   NAND4_X1 i_848 (.A1(in2[24]), .A2(in2[23]), .A3(in1[22]), .A4(in1[21]), 
      .ZN(n_832));
   AOI22_X1 i_849 (.A1(in2[24]), .A2(in1[21]), .B1(in2[23]), .B2(in1[22]), 
      .ZN(n_833));
   NAND2_X1 i_850 (.A1(in2[25]), .A2(in1[20]), .ZN(n_834));
   OAI21_X1 i_851 (.A(n_832), .B1(n_833), .B2(n_834), .ZN(n_454));
   NAND4_X1 i_852 (.A1(in1[25]), .A2(in1[24]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_835));
   AOI22_X1 i_853 (.A1(in1[24]), .A2(in2[21]), .B1(in1[25]), .B2(in2[20]), 
      .ZN(n_836));
   NAND2_X1 i_854 (.A1(in1[23]), .A2(in2[22]), .ZN(n_837));
   OAI21_X1 i_855 (.A(n_835), .B1(n_836), .B2(n_837), .ZN(n_455));
   NAND4_X1 i_856 (.A1(in1[28]), .A2(in1[27]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_838));
   AOI22_X1 i_857 (.A1(in1[27]), .A2(in2[18]), .B1(in1[28]), .B2(in2[17]), 
      .ZN(n_839));
   NAND2_X1 i_858 (.A1(in1[26]), .A2(in2[19]), .ZN(n_840));
   OAI21_X1 i_859 (.A(n_838), .B1(n_839), .B2(n_840), .ZN(n_456));
   INV_X1 i_860 (.A(n_826), .ZN(n_841));
   NAND2_X1 i_861 (.A1(n_841), .A2(n_825), .ZN(n_842));
   XOR2_X1 i_862 (.A(n_842), .B(n_827), .Z(n_457));
   INV_X1 i_863 (.A(n_829), .ZN(n_843));
   NAND2_X1 i_864 (.A1(n_843), .A2(n_828), .ZN(n_844));
   XOR2_X1 i_865 (.A(n_844), .B(n_830), .Z(n_458));
   INV_X1 i_866 (.A(n_833), .ZN(n_845));
   NAND2_X1 i_867 (.A1(n_845), .A2(n_832), .ZN(n_846));
   XOR2_X1 i_868 (.A(n_846), .B(n_834), .Z(n_459));
   INV_X1 i_869 (.A(n_836), .ZN(n_847));
   NAND2_X1 i_870 (.A1(n_847), .A2(n_835), .ZN(n_848));
   XOR2_X1 i_871 (.A(n_848), .B(n_837), .Z(n_460));
   INV_X1 i_872 (.A(n_839), .ZN(n_849));
   NAND2_X1 i_873 (.A1(n_849), .A2(n_838), .ZN(n_850));
   XOR2_X1 i_874 (.A(n_850), .B(n_840), .Z(n_461));
   NAND2_X1 i_875 (.A1(n_789), .A2(n_791), .ZN(n_851));
   XOR2_X1 i_876 (.A(n_851), .B(n_793), .Z(n_462));
   NAND4_X1 i_877 (.A1(in2[30]), .A2(in2[29]), .A3(in1[14]), .A4(in1[15]), 
      .ZN(n_852));
   AOI22_X1 i_878 (.A1(in2[30]), .A2(in1[14]), .B1(in2[29]), .B2(in1[15]), 
      .ZN(n_853));
   AND2_X1 i_879 (.A1(in2[31]), .A2(in1[13]), .ZN(n_854));
   OAI21_X1 i_880 (.A(n_852), .B1(n_853), .B2(n_854), .ZN(n_463));
   NAND4_X1 i_881 (.A1(in2[27]), .A2(in2[26]), .A3(in1[17]), .A4(in1[18]), 
      .ZN(n_855));
   AOI22_X1 i_882 (.A1(in2[27]), .A2(in1[17]), .B1(in2[26]), .B2(in1[18]), 
      .ZN(n_856));
   NAND2_X1 i_883 (.A1(in2[28]), .A2(in1[16]), .ZN(n_857));
   OAI21_X1 i_884 (.A(n_855), .B1(n_856), .B2(n_857), .ZN(n_464));
   NAND4_X1 i_885 (.A1(in2[24]), .A2(in2[23]), .A3(in1[20]), .A4(in1[21]), 
      .ZN(n_858));
   AOI22_X1 i_886 (.A1(in2[24]), .A2(in1[20]), .B1(in2[23]), .B2(in1[21]), 
      .ZN(n_859));
   NAND2_X1 i_887 (.A1(in2[25]), .A2(in1[19]), .ZN(n_860));
   OAI21_X1 i_888 (.A(n_858), .B1(n_859), .B2(n_860), .ZN(n_465));
   NAND4_X1 i_889 (.A1(in1[23]), .A2(in1[24]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_861));
   AOI22_X1 i_890 (.A1(in1[23]), .A2(in2[21]), .B1(in1[24]), .B2(in2[20]), 
      .ZN(n_862));
   NAND2_X1 i_891 (.A1(in1[22]), .A2(in2[22]), .ZN(n_863));
   OAI21_X1 i_892 (.A(n_861), .B1(n_862), .B2(n_863), .ZN(n_466));
   NAND4_X1 i_893 (.A1(in1[26]), .A2(in1[27]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_864));
   AOI22_X1 i_894 (.A1(in1[26]), .A2(in2[18]), .B1(in1[27]), .B2(in2[17]), 
      .ZN(n_865));
   NAND2_X1 i_895 (.A1(in1[25]), .A2(in2[19]), .ZN(n_866));
   OAI21_X1 i_896 (.A(n_864), .B1(n_865), .B2(n_866), .ZN(n_467));
   NAND4_X1 i_897 (.A1(in1[29]), .A2(in1[30]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_867));
   AOI22_X1 i_898 (.A1(in1[29]), .A2(in2[15]), .B1(in1[30]), .B2(in2[14]), 
      .ZN(n_868));
   NAND2_X1 i_899 (.A1(in1[28]), .A2(in2[16]), .ZN(n_869));
   OAI21_X1 i_900 (.A(n_867), .B1(n_868), .B2(n_869), .ZN(n_468));
   INV_X1 i_901 (.A(n_853), .ZN(n_870));
   NAND2_X1 i_902 (.A1(n_870), .A2(n_852), .ZN(n_871));
   XOR2_X1 i_903 (.A(n_871), .B(n_854), .Z(n_469));
   INV_X1 i_904 (.A(n_856), .ZN(n_872));
   NAND2_X1 i_905 (.A1(n_872), .A2(n_855), .ZN(n_873));
   XOR2_X1 i_906 (.A(n_873), .B(n_857), .Z(n_470));
   INV_X1 i_907 (.A(n_859), .ZN(n_874));
   NAND2_X1 i_908 (.A1(n_874), .A2(n_858), .ZN(n_875));
   XOR2_X1 i_909 (.A(n_875), .B(n_860), .Z(n_471));
   INV_X1 i_910 (.A(n_862), .ZN(n_876));
   NAND2_X1 i_911 (.A1(n_876), .A2(n_861), .ZN(n_877));
   XOR2_X1 i_912 (.A(n_877), .B(n_863), .Z(n_472));
   INV_X1 i_913 (.A(n_865), .ZN(n_878));
   NAND2_X1 i_914 (.A1(n_878), .A2(n_864), .ZN(n_879));
   XOR2_X1 i_915 (.A(n_879), .B(n_866), .Z(n_473));
   INV_X1 i_916 (.A(n_868), .ZN(n_880));
   NAND2_X1 i_917 (.A1(n_880), .A2(n_867), .ZN(n_881));
   XOR2_X1 i_918 (.A(n_881), .B(n_869), .Z(n_474));
   NAND4_X1 i_919 (.A1(in2[30]), .A2(in2[29]), .A3(in1[14]), .A4(in1[13]), 
      .ZN(n_894));
   AOI22_X1 i_920 (.A1(in2[30]), .A2(in1[13]), .B1(in2[29]), .B2(in1[14]), 
      .ZN(n_895));
   AND2_X1 i_921 (.A1(in2[31]), .A2(in1[12]), .ZN(n_896));
   OAI21_X1 i_922 (.A(n_894), .B1(n_895), .B2(n_896), .ZN(n_476));
   NAND4_X1 i_923 (.A1(in2[27]), .A2(in2[26]), .A3(in1[17]), .A4(in1[16]), 
      .ZN(n_897));
   AOI22_X1 i_924 (.A1(in2[27]), .A2(in1[16]), .B1(in2[26]), .B2(in1[17]), 
      .ZN(n_898));
   NAND2_X1 i_925 (.A1(in2[28]), .A2(in1[15]), .ZN(n_899));
   OAI21_X1 i_926 (.A(n_897), .B1(n_898), .B2(n_899), .ZN(n_477));
   NAND4_X1 i_927 (.A1(in2[24]), .A2(in2[23]), .A3(in1[20]), .A4(in1[19]), 
      .ZN(n_900));
   AOI22_X1 i_928 (.A1(in2[24]), .A2(in1[19]), .B1(in2[23]), .B2(in1[20]), 
      .ZN(n_901));
   NAND2_X1 i_929 (.A1(in2[25]), .A2(in1[18]), .ZN(n_902));
   OAI21_X1 i_930 (.A(n_900), .B1(n_901), .B2(n_902), .ZN(n_478));
   NAND4_X1 i_931 (.A1(in1[23]), .A2(in1[22]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_903));
   AOI22_X1 i_932 (.A1(in1[22]), .A2(in2[21]), .B1(in1[23]), .B2(in2[20]), 
      .ZN(n_904));
   NAND2_X1 i_933 (.A1(in2[22]), .A2(in1[21]), .ZN(n_905));
   OAI21_X1 i_934 (.A(n_903), .B1(n_904), .B2(n_905), .ZN(n_479));
   NAND4_X1 i_935 (.A1(in1[26]), .A2(in1[25]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_906));
   AOI22_X1 i_936 (.A1(in1[25]), .A2(in2[18]), .B1(in1[26]), .B2(in2[17]), 
      .ZN(n_907));
   NAND2_X1 i_937 (.A1(in1[24]), .A2(in2[19]), .ZN(n_908));
   OAI21_X1 i_938 (.A(n_906), .B1(n_907), .B2(n_908), .ZN(n_480));
   NOR2_X1 i_939 (.A1(n_1580), .A2(n_790), .ZN(n_909));
   NAND3_X1 i_940 (.A1(n_909), .A2(in1[29]), .A3(in2[14]), .ZN(n_910));
   AOI21_X1 i_941 (.A(n_909), .B1(in1[29]), .B2(in2[14]), .ZN(n_911));
   NAND2_X1 i_942 (.A1(in1[27]), .A2(in2[16]), .ZN(n_912));
   OAI21_X1 i_943 (.A(n_910), .B1(n_911), .B2(n_912), .ZN(n_481));
   NAND2_X1 i_944 (.A1(in1[31]), .A2(in2[13]), .ZN(n_482));
   INV_X1 i_945 (.A(n_895), .ZN(n_913));
   NAND2_X1 i_946 (.A1(n_913), .A2(n_894), .ZN(n_914));
   XOR2_X1 i_947 (.A(n_914), .B(n_896), .Z(n_483));
   INV_X1 i_948 (.A(n_898), .ZN(n_915));
   NAND2_X1 i_949 (.A1(n_915), .A2(n_897), .ZN(n_916));
   XOR2_X1 i_950 (.A(n_916), .B(n_899), .Z(n_484));
   INV_X1 i_951 (.A(n_901), .ZN(n_917));
   NAND2_X1 i_952 (.A1(n_917), .A2(n_900), .ZN(n_918));
   XOR2_X1 i_953 (.A(n_918), .B(n_902), .Z(n_485));
   INV_X1 i_954 (.A(n_904), .ZN(n_919));
   NAND2_X1 i_955 (.A1(n_919), .A2(n_903), .ZN(n_920));
   XOR2_X1 i_956 (.A(n_920), .B(n_905), .Z(n_486));
   INV_X1 i_957 (.A(n_907), .ZN(n_921));
   NAND2_X1 i_958 (.A1(n_921), .A2(n_906), .ZN(n_922));
   XOR2_X1 i_959 (.A(n_922), .B(n_908), .Z(n_487));
   INV_X1 i_960 (.A(n_911), .ZN(n_923));
   NAND2_X1 i_961 (.A1(n_910), .A2(n_923), .ZN(n_924));
   XOR2_X1 i_962 (.A(n_924), .B(n_912), .Z(n_488));
   XNOR2_X1 i_963 (.A(n_2086), .B(n_2092), .ZN(n_489));
   NAND4_X1 i_964 (.A1(in2[30]), .A2(in2[29]), .A3(in1[13]), .A4(in1[12]), 
      .ZN(n_925));
   AOI22_X1 i_965 (.A1(in2[30]), .A2(in1[12]), .B1(in2[29]), .B2(in1[13]), 
      .ZN(n_926));
   AND2_X1 i_966 (.A1(in2[31]), .A2(in1[11]), .ZN(n_928));
   OAI21_X1 i_967 (.A(n_925), .B1(n_926), .B2(n_928), .ZN(n_490));
   NAND4_X1 i_968 (.A1(in2[27]), .A2(in2[26]), .A3(in1[16]), .A4(in1[15]), 
      .ZN(n_929));
   AOI22_X1 i_969 (.A1(in2[27]), .A2(in1[15]), .B1(in2[26]), .B2(in1[16]), 
      .ZN(n_930));
   NAND2_X1 i_970 (.A1(in2[28]), .A2(in1[14]), .ZN(n_931));
   OAI21_X1 i_971 (.A(n_929), .B1(n_930), .B2(n_931), .ZN(n_491));
   NAND4_X1 i_972 (.A1(in2[24]), .A2(in2[23]), .A3(in1[19]), .A4(in1[18]), 
      .ZN(n_932));
   AOI22_X1 i_973 (.A1(in2[24]), .A2(in1[18]), .B1(in2[23]), .B2(in1[19]), 
      .ZN(n_933));
   NAND2_X1 i_974 (.A1(in2[25]), .A2(in1[17]), .ZN(n_934));
   OAI21_X1 i_975 (.A(n_932), .B1(n_933), .B2(n_934), .ZN(n_492));
   NAND4_X1 i_976 (.A1(in1[22]), .A2(in1[21]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_935));
   AOI22_X1 i_977 (.A1(in1[21]), .A2(in2[21]), .B1(in1[22]), .B2(in2[20]), 
      .ZN(n_936));
   NAND2_X1 i_978 (.A1(in2[22]), .A2(in1[20]), .ZN(n_937));
   OAI21_X1 i_979 (.A(n_935), .B1(n_936), .B2(n_937), .ZN(n_493));
   NAND4_X1 i_980 (.A1(in1[25]), .A2(in1[24]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_938));
   AOI22_X1 i_981 (.A1(in1[24]), .A2(in2[18]), .B1(in1[25]), .B2(in2[17]), 
      .ZN(n_939));
   NAND2_X1 i_982 (.A1(in1[23]), .A2(in2[19]), .ZN(n_940));
   OAI21_X1 i_983 (.A(n_938), .B1(n_939), .B2(n_940), .ZN(n_494));
   NAND4_X1 i_984 (.A1(in1[28]), .A2(in1[27]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_941));
   AOI22_X1 i_985 (.A1(in1[27]), .A2(in2[15]), .B1(in1[28]), .B2(in2[14]), 
      .ZN(n_942));
   NAND2_X1 i_986 (.A1(in1[26]), .A2(in2[16]), .ZN(n_943));
   OAI21_X1 i_987 (.A(n_941), .B1(n_942), .B2(n_943), .ZN(n_495));
   INV_X1 i_988 (.A(n_926), .ZN(n_944));
   NAND2_X1 i_989 (.A1(n_944), .A2(n_925), .ZN(n_945));
   XOR2_X1 i_990 (.A(n_945), .B(n_928), .Z(n_496));
   INV_X1 i_991 (.A(n_930), .ZN(n_946));
   NAND2_X1 i_992 (.A1(n_946), .A2(n_929), .ZN(n_947));
   XOR2_X1 i_993 (.A(n_947), .B(n_931), .Z(n_497));
   INV_X1 i_994 (.A(n_933), .ZN(n_948));
   NAND2_X1 i_995 (.A1(n_948), .A2(n_932), .ZN(n_949));
   XOR2_X1 i_996 (.A(n_949), .B(n_934), .Z(n_498));
   INV_X1 i_997 (.A(n_936), .ZN(n_950));
   NAND2_X1 i_998 (.A1(n_950), .A2(n_935), .ZN(n_951));
   XOR2_X1 i_999 (.A(n_951), .B(n_937), .Z(n_499));
   INV_X1 i_1000 (.A(n_939), .ZN(n_952));
   NAND2_X1 i_1001 (.A1(n_952), .A2(n_938), .ZN(n_953));
   XOR2_X1 i_1002 (.A(n_953), .B(n_940), .Z(n_500));
   INV_X1 i_1003 (.A(n_942), .ZN(n_954));
   NAND2_X1 i_1004 (.A1(n_954), .A2(n_941), .ZN(n_955));
   XOR2_X1 i_1005 (.A(n_955), .B(n_943), .Z(n_501));
   NAND2_X1 i_1006 (.A1(n_2258), .A2(n_2257), .ZN(n_956));
   XOR2_X1 i_1007 (.A(n_956), .B(n_2093), .Z(n_502));
   NAND4_X1 i_1008 (.A1(in2[30]), .A2(in2[29]), .A3(in1[11]), .A4(in1[12]), 
      .ZN(n_957));
   AOI22_X1 i_1009 (.A1(in2[30]), .A2(in1[11]), .B1(in2[29]), .B2(in1[12]), 
      .ZN(n_958));
   AND2_X1 i_1010 (.A1(in2[31]), .A2(in1[10]), .ZN(n_959));
   OAI21_X1 i_1011 (.A(n_957), .B1(n_958), .B2(n_959), .ZN(n_391));
   NAND4_X1 i_1012 (.A1(in2[27]), .A2(in2[26]), .A3(in1[14]), .A4(in1[15]), 
      .ZN(n_960));
   AOI22_X1 i_1013 (.A1(in2[27]), .A2(in1[14]), .B1(in2[26]), .B2(in1[15]), 
      .ZN(n_961));
   NAND2_X1 i_1014 (.A1(in2[28]), .A2(in1[13]), .ZN(n_962));
   OAI21_X1 i_1015 (.A(n_960), .B1(n_961), .B2(n_962), .ZN(n_503));
   NAND4_X1 i_1016 (.A1(in2[24]), .A2(in2[23]), .A3(in1[17]), .A4(in1[18]), 
      .ZN(n_963));
   AOI22_X1 i_1017 (.A1(in2[24]), .A2(in1[17]), .B1(in2[23]), .B2(in1[18]), 
      .ZN(n_964));
   NAND2_X1 i_1018 (.A1(in2[25]), .A2(in1[16]), .ZN(n_965));
   OAI21_X1 i_1019 (.A(n_963), .B1(n_964), .B2(n_965), .ZN(n_504));
   NAND4_X1 i_1020 (.A1(in1[20]), .A2(in1[21]), .A3(in2[21]), .A4(in2[20]), 
      .ZN(n_966));
   AOI22_X1 i_1021 (.A1(in1[20]), .A2(in2[21]), .B1(in1[21]), .B2(in2[20]), 
      .ZN(n_967));
   NAND2_X1 i_1022 (.A1(in2[22]), .A2(in1[19]), .ZN(n_968));
   OAI21_X1 i_1023 (.A(n_966), .B1(n_967), .B2(n_968), .ZN(n_505));
   NAND4_X1 i_1024 (.A1(in1[23]), .A2(in1[24]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_969));
   AOI22_X1 i_1025 (.A1(in1[23]), .A2(in2[18]), .B1(in1[24]), .B2(in2[17]), 
      .ZN(n_970));
   NAND2_X1 i_1026 (.A1(in1[22]), .A2(in2[19]), .ZN(n_971));
   OAI21_X1 i_1027 (.A(n_969), .B1(n_970), .B2(n_971), .ZN(n_506));
   NAND4_X1 i_1028 (.A1(in1[26]), .A2(in1[27]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_972));
   AOI22_X1 i_1029 (.A1(in1[26]), .A2(in2[15]), .B1(in1[27]), .B2(in2[14]), 
      .ZN(n_973));
   NAND2_X1 i_1030 (.A1(in1[25]), .A2(in2[16]), .ZN(n_974));
   OAI21_X1 i_1031 (.A(n_972), .B1(n_973), .B2(n_974), .ZN(n_507));
   NAND4_X1 i_1032 (.A1(in1[29]), .A2(in1[30]), .A3(in2[12]), .A4(in2[11]), 
      .ZN(n_975));
   AOI22_X1 i_1033 (.A1(in1[29]), .A2(in2[12]), .B1(in1[30]), .B2(in2[11]), 
      .ZN(n_976));
   NAND2_X1 i_1034 (.A1(in1[28]), .A2(in2[13]), .ZN(n_977));
   OAI21_X1 i_1035 (.A(n_975), .B1(n_976), .B2(n_977), .ZN(n_508));
   INV_X1 i_1036 (.A(n_958), .ZN(n_978));
   NAND2_X1 i_1037 (.A1(n_978), .A2(n_957), .ZN(n_979));
   XOR2_X1 i_1038 (.A(n_979), .B(n_959), .Z(n_394));
   INV_X1 i_1039 (.A(n_961), .ZN(n_980));
   NAND2_X1 i_1040 (.A1(n_980), .A2(n_960), .ZN(n_981));
   XOR2_X1 i_1041 (.A(n_981), .B(n_962), .Z(n_509));
   INV_X1 i_1042 (.A(n_964), .ZN(n_982));
   NAND2_X1 i_1043 (.A1(n_982), .A2(n_963), .ZN(n_983));
   XOR2_X1 i_1044 (.A(n_983), .B(n_965), .Z(n_510));
   INV_X1 i_1045 (.A(n_967), .ZN(n_984));
   NAND2_X1 i_1046 (.A1(n_984), .A2(n_966), .ZN(n_985));
   XOR2_X1 i_1047 (.A(n_985), .B(n_968), .Z(n_511));
   INV_X1 i_1048 (.A(n_970), .ZN(n_986));
   NAND2_X1 i_1049 (.A1(n_986), .A2(n_969), .ZN(n_987));
   XOR2_X1 i_1050 (.A(n_987), .B(n_971), .Z(n_512));
   INV_X1 i_1051 (.A(n_973), .ZN(n_988));
   NAND2_X1 i_1052 (.A1(n_988), .A2(n_972), .ZN(n_989));
   XOR2_X1 i_1053 (.A(n_989), .B(n_974), .Z(n_513));
   INV_X1 i_1054 (.A(n_976), .ZN(n_990));
   NAND2_X1 i_1055 (.A1(n_990), .A2(n_975), .ZN(n_992));
   XOR2_X1 i_1056 (.A(n_992), .B(n_977), .Z(n_514));
   AND2_X1 i_1057 (.A1(in1[30]), .A2(in2[10]), .ZN(n_993));
   INV_X1 i_1058 (.A(in2[8]), .ZN(n_994));
   OAI211_X1 i_1059 (.A(in1[30]), .B(in2[9]), .C1(n_1384), .C2(n_994), .ZN(n_995));
   INV_X1 i_1060 (.A(in2[9]), .ZN(n_996));
   OAI211_X1 i_1061 (.A(in1[31]), .B(in2[8]), .C1(n_1383), .C2(n_996), .ZN(n_997));
   INV_X1 i_1062 (.A(n_997), .ZN(n_998));
   NAND2_X1 i_1063 (.A1(in1[29]), .A2(in2[10]), .ZN(n_999));
   OAI21_X1 i_1064 (.A(n_995), .B1(n_998), .B2(n_999), .ZN(n_1000));
   NOR2_X1 i_1065 (.A1(n_1384), .A2(n_996), .ZN(n_1001));
   XOR2_X1 i_1066 (.A(n_993), .B(n_1001), .Z(n_1002));
   OAI21_X1 i_1067 (.A(n_993), .B1(n_1000), .B2(n_1002), .ZN(n_1003));
   INV_X1 i_1068 (.A(n_1000), .ZN(n_1004));
   OAI21_X1 i_1069 (.A(n_1003), .B1(n_1004), .B2(n_1001), .ZN(n_395));
   NAND4_X1 i_1070 (.A1(in2[30]), .A2(in2[29]), .A3(in1[11]), .A4(in1[10]), 
      .ZN(n_1005));
   AOI22_X1 i_1071 (.A1(in2[30]), .A2(in1[10]), .B1(in2[29]), .B2(in1[11]), 
      .ZN(n_1006));
   AND2_X1 i_1072 (.A1(in2[31]), .A2(in1[9]), .ZN(n_1007));
   OAI21_X1 i_1073 (.A(n_1005), .B1(n_1006), .B2(n_1007), .ZN(n_3697));
   NAND4_X1 i_1074 (.A1(in2[27]), .A2(in2[26]), .A3(in1[14]), .A4(in1[13]), 
      .ZN(n_1008));
   AOI22_X1 i_1075 (.A1(in2[27]), .A2(in1[13]), .B1(in2[26]), .B2(in1[14]), 
      .ZN(n_1009));
   NAND2_X1 i_1076 (.A1(in2[28]), .A2(in1[12]), .ZN(n_1010));
   OAI21_X1 i_1077 (.A(n_1008), .B1(n_1009), .B2(n_1010), .ZN(n_3706));
   NAND4_X1 i_1078 (.A1(in2[24]), .A2(in2[23]), .A3(in1[17]), .A4(in1[16]), 
      .ZN(n_1011));
   AOI22_X1 i_1079 (.A1(in2[24]), .A2(in1[16]), .B1(in2[23]), .B2(in1[17]), 
      .ZN(n_1012));
   NAND2_X1 i_1080 (.A1(in2[25]), .A2(in1[15]), .ZN(n_1013));
   OAI21_X1 i_1081 (.A(n_1011), .B1(n_1012), .B2(n_1013), .ZN(n_3713));
   NAND4_X1 i_1082 (.A1(in1[20]), .A2(in2[21]), .A3(in2[20]), .A4(in1[19]), 
      .ZN(n_1014));
   AOI22_X1 i_1083 (.A1(in2[21]), .A2(in1[19]), .B1(in1[20]), .B2(in2[20]), 
      .ZN(n_1015));
   NAND2_X1 i_1084 (.A1(in2[22]), .A2(in1[18]), .ZN(n_1016));
   OAI21_X1 i_1085 (.A(n_1014), .B1(n_1015), .B2(n_1016), .ZN(n_3720));
   NAND4_X1 i_1086 (.A1(in1[23]), .A2(in1[22]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_1017));
   AOI22_X1 i_1087 (.A1(in1[22]), .A2(in2[18]), .B1(in1[23]), .B2(in2[17]), 
      .ZN(n_1018));
   NAND2_X1 i_1088 (.A1(in1[21]), .A2(in2[19]), .ZN(n_1019));
   OAI21_X1 i_1089 (.A(n_1017), .B1(n_1018), .B2(n_1019), .ZN(n_3727));
   NAND4_X1 i_1090 (.A1(in1[26]), .A2(in1[25]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_1020));
   AOI22_X1 i_1091 (.A1(in1[25]), .A2(in2[15]), .B1(in1[26]), .B2(in2[14]), 
      .ZN(n_1021));
   NAND2_X1 i_1092 (.A1(in1[24]), .A2(in2[16]), .ZN(n_1023));
   OAI21_X1 i_1093 (.A(n_1020), .B1(n_1021), .B2(n_1023), .ZN(n_3734));
   NOR2_X1 i_1094 (.A1(n_1580), .A2(n_2262), .ZN(n_1024));
   NAND3_X1 i_1095 (.A1(n_1024), .A2(in1[29]), .A3(in2[11]), .ZN(n_1025));
   AOI21_X1 i_1096 (.A(n_1024), .B1(in1[29]), .B2(in2[11]), .ZN(n_1026));
   NAND2_X1 i_1097 (.A1(in1[27]), .A2(in2[13]), .ZN(n_1027));
   OAI21_X1 i_1098 (.A(n_1025), .B1(n_1026), .B2(n_1027), .ZN(n_396));
   NAND2_X1 i_1099 (.A1(in1[31]), .A2(in2[10]), .ZN(n_515));
   INV_X1 i_1100 (.A(n_1006), .ZN(n_1028));
   NAND2_X1 i_1101 (.A1(n_1028), .A2(n_1005), .ZN(n_1031));
   XOR2_X1 i_1102 (.A(n_1031), .B(n_1007), .Z(n_3696));
   INV_X1 i_1103 (.A(n_1009), .ZN(n_1032));
   NAND2_X1 i_1104 (.A1(n_1032), .A2(n_1008), .ZN(n_1033));
   XOR2_X1 i_1105 (.A(n_1033), .B(n_1010), .Z(n_3705));
   INV_X1 i_1106 (.A(n_1012), .ZN(n_1035));
   NAND2_X1 i_1107 (.A1(n_1035), .A2(n_1011), .ZN(n_1036));
   XOR2_X1 i_1108 (.A(n_1036), .B(n_1013), .Z(n_3712));
   INV_X1 i_1109 (.A(n_1015), .ZN(n_1037));
   NAND2_X1 i_1110 (.A1(n_1037), .A2(n_1014), .ZN(n_1038));
   XOR2_X1 i_1111 (.A(n_1038), .B(n_1016), .Z(n_3719));
   INV_X1 i_1112 (.A(n_1018), .ZN(n_1041));
   NAND2_X1 i_1113 (.A1(n_1041), .A2(n_1017), .ZN(n_1042));
   XOR2_X1 i_1114 (.A(n_1042), .B(n_1019), .Z(n_3726));
   INV_X1 i_1115 (.A(n_1021), .ZN(n_1043));
   NAND2_X1 i_1116 (.A1(n_1043), .A2(n_1020), .ZN(n_1044));
   XOR2_X1 i_1117 (.A(n_1044), .B(n_1023), .Z(n_3733));
   INV_X1 i_1118 (.A(n_1026), .ZN(n_1047));
   NAND2_X1 i_1119 (.A1(n_1025), .A2(n_1047), .ZN(n_1048));
   XOR2_X1 i_1120 (.A(n_1048), .B(n_1027), .Z(n_397));
   XNOR2_X1 i_1121 (.A(n_1002), .B(n_1000), .ZN(n_398));
   OAI21_X1 i_1122 (.A(n_2077), .B1(n_2078), .B2(n_2076), .ZN(n_3609));
   NAND4_X1 i_1123 (.A1(in2[27]), .A2(in2[26]), .A3(in1[13]), .A4(in1[12]), 
      .ZN(n_1054));
   AOI22_X1 i_1124 (.A1(in2[27]), .A2(in1[12]), .B1(in2[26]), .B2(in1[13]), 
      .ZN(n_1055));
   NAND2_X1 i_1125 (.A1(in2[28]), .A2(in1[11]), .ZN(n_1057));
   OAI21_X1 i_1126 (.A(n_1054), .B1(n_1055), .B2(n_1057), .ZN(n_3618));
   NAND4_X1 i_1127 (.A1(in2[24]), .A2(in2[23]), .A3(in1[16]), .A4(in1[15]), 
      .ZN(n_1058));
   AOI22_X1 i_1128 (.A1(in2[24]), .A2(in1[15]), .B1(in2[23]), .B2(in1[16]), 
      .ZN(n_1059));
   NAND2_X1 i_1129 (.A1(in2[25]), .A2(in1[14]), .ZN(n_1060));
   OAI21_X1 i_1130 (.A(n_1058), .B1(n_1059), .B2(n_1060), .ZN(n_3625));
   NAND4_X1 i_1131 (.A1(in2[21]), .A2(in2[20]), .A3(in1[19]), .A4(in1[18]), 
      .ZN(n_1061));
   AOI22_X1 i_1132 (.A1(in2[21]), .A2(in1[18]), .B1(in2[20]), .B2(in1[19]), 
      .ZN(n_1062));
   NAND2_X1 i_1133 (.A1(in2[22]), .A2(in1[17]), .ZN(n_1064));
   OAI21_X1 i_1134 (.A(n_1061), .B1(n_1062), .B2(n_1064), .ZN(n_3632));
   NAND4_X1 i_1135 (.A1(in1[22]), .A2(in1[21]), .A3(in2[18]), .A4(in2[17]), 
      .ZN(n_1065));
   AOI22_X1 i_1136 (.A1(in1[21]), .A2(in2[18]), .B1(in1[22]), .B2(in2[17]), 
      .ZN(n_1066));
   NAND2_X1 i_1137 (.A1(in1[20]), .A2(in2[19]), .ZN(n_1067));
   OAI21_X1 i_1138 (.A(n_1065), .B1(n_1066), .B2(n_1067), .ZN(n_3639));
   NAND4_X1 i_1139 (.A1(in1[25]), .A2(in1[24]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_1072));
   AOI22_X1 i_1140 (.A1(in1[24]), .A2(in2[15]), .B1(in1[25]), .B2(in2[14]), 
      .ZN(n_1073));
   NAND2_X1 i_1141 (.A1(in1[23]), .A2(in2[16]), .ZN(n_1076));
   OAI21_X1 i_1142 (.A(n_1072), .B1(n_1073), .B2(n_1076), .ZN(n_3646));
   NAND4_X1 i_1143 (.A1(in1[28]), .A2(in1[27]), .A3(in2[12]), .A4(in2[11]), 
      .ZN(n_1077));
   AOI22_X1 i_1144 (.A1(in1[27]), .A2(in2[12]), .B1(in1[28]), .B2(in2[11]), 
      .ZN(n_1078));
   NAND2_X1 i_1145 (.A1(in1[26]), .A2(in2[13]), .ZN(n_1079));
   OAI21_X1 i_1146 (.A(n_1077), .B1(n_1078), .B2(n_1079), .ZN(n_3653));
   INV_X1 i_1147 (.A(n_1055), .ZN(n_1083));
   NAND2_X1 i_1148 (.A1(n_1083), .A2(n_1054), .ZN(n_1084));
   XOR2_X1 i_1149 (.A(n_1084), .B(n_1057), .Z(n_3617));
   INV_X1 i_1150 (.A(n_1059), .ZN(n_1085));
   NAND2_X1 i_1151 (.A1(n_1085), .A2(n_1058), .ZN(n_1086));
   XOR2_X1 i_1152 (.A(n_1086), .B(n_1060), .Z(n_3624));
   INV_X1 i_1153 (.A(n_1062), .ZN(n_1087));
   NAND2_X1 i_1154 (.A1(n_1087), .A2(n_1061), .ZN(n_1090));
   XOR2_X1 i_1155 (.A(n_1090), .B(n_1064), .Z(n_3631));
   INV_X1 i_1156 (.A(n_1066), .ZN(n_1091));
   NAND2_X1 i_1157 (.A1(n_1091), .A2(n_1065), .ZN(n_1092));
   XOR2_X1 i_1158 (.A(n_1092), .B(n_1067), .Z(n_3638));
   INV_X1 i_1159 (.A(n_1073), .ZN(n_1093));
   NAND2_X1 i_1160 (.A1(n_1093), .A2(n_1072), .ZN(n_1098));
   XOR2_X1 i_1161 (.A(n_1098), .B(n_1076), .Z(n_3645));
   INV_X1 i_1162 (.A(n_1078), .ZN(n_1099));
   NAND2_X1 i_1163 (.A1(n_1099), .A2(n_1077), .ZN(n_1102));
   XOR2_X1 i_1164 (.A(n_1102), .B(n_1079), .Z(n_3652));
   NAND2_X1 i_1165 (.A1(n_995), .A2(n_997), .ZN(n_1103));
   XOR2_X1 i_1166 (.A(n_1103), .B(n_999), .Z(n_3658));
   NAND3_X1 i_1167 (.A1(n_1938), .A2(in2[24]), .A3(in1[15]), .ZN(n_1116));
   AOI22_X1 i_1168 (.A1(in2[24]), .A2(in1[14]), .B1(in2[23]), .B2(in1[15]), 
      .ZN(n_1117));
   NAND2_X1 i_1169 (.A1(in2[25]), .A2(in1[13]), .ZN(n_1118));
   OAI21_X1 i_1170 (.A(n_1116), .B1(n_1117), .B2(n_1118), .ZN(n_3536));
   NAND4_X1 i_1171 (.A1(in2[21]), .A2(in2[20]), .A3(in1[17]), .A4(in1[18]), 
      .ZN(n_1119));
   AOI22_X1 i_1172 (.A1(in2[21]), .A2(in1[17]), .B1(in2[20]), .B2(in1[18]), 
      .ZN(n_1126));
   NAND2_X1 i_1175 (.A1(in2[22]), .A2(in1[16]), .ZN(n_1127));
   OAI21_X1 i_1176 (.A(n_1119), .B1(n_1126), .B2(n_1127), .ZN(n_3543));
   AND2_X1 i_1177 (.A1(in1[20]), .A2(in2[17]), .ZN(n_1130));
   NAND3_X1 i_1178 (.A1(n_1130), .A2(in1[21]), .A3(in2[18]), .ZN(n_1131));
   AOI22_X1 i_1179 (.A1(in1[20]), .A2(in2[18]), .B1(in1[21]), .B2(in2[17]), 
      .ZN(n_1132));
   NAND2_X1 i_1180 (.A1(in1[19]), .A2(in2[19]), .ZN(n_1133));
   OAI21_X1 i_1181 (.A(n_1131), .B1(n_1132), .B2(n_1133), .ZN(n_3550));
   NAND4_X1 i_1182 (.A1(in1[23]), .A2(in1[24]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_1134));
   AOI22_X1 i_1183 (.A1(in1[23]), .A2(in2[15]), .B1(in1[24]), .B2(in2[14]), 
      .ZN(n_1136));
   NAND2_X1 i_1184 (.A1(in1[22]), .A2(in2[16]), .ZN(n_1137));
   OAI21_X1 i_1185 (.A(n_1134), .B1(n_1136), .B2(n_1137), .ZN(n_3557));
   AND2_X1 i_1186 (.A1(in1[26]), .A2(in2[11]), .ZN(n_1138));
   NAND3_X1 i_1187 (.A1(n_1138), .A2(in1[27]), .A3(in2[12]), .ZN(n_1139));
   AOI22_X1 i_1188 (.A1(in1[26]), .A2(in2[12]), .B1(in1[27]), .B2(in2[11]), 
      .ZN(n_1140));
   NAND2_X1 i_1189 (.A1(in1[25]), .A2(in2[13]), .ZN(n_1141));
   OAI21_X1 i_1190 (.A(n_1139), .B1(n_1140), .B2(n_1141), .ZN(n_3564));
   NOR2_X1 i_1191 (.A1(n_1382), .A2(n_994), .ZN(n_1143));
   NAND3_X1 i_1192 (.A1(n_1143), .A2(in1[30]), .A3(in2[9]), .ZN(n_1144));
   AOI22_X1 i_1193 (.A1(in1[29]), .A2(in2[9]), .B1(in1[30]), .B2(in2[8]), 
      .ZN(n_1145));
   NAND2_X1 i_1194 (.A1(in1[28]), .A2(in2[10]), .ZN(n_1146));
   OAI21_X1 i_1195 (.A(n_1144), .B1(n_1145), .B2(n_1146), .ZN(n_3571));
   INV_X1 i_1196 (.A(n_1940), .ZN(n_1155));
   NAND2_X1 i_1197 (.A1(n_1155), .A2(n_1941), .ZN(n_1156));
   XOR2_X1 i_1198 (.A(n_1156), .B(n_1939), .Z(n_3519));
   INV_X1 i_1199 (.A(n_1945), .ZN(n_1159));
   NAND2_X1 i_1200 (.A1(n_1946), .A2(n_1159), .ZN(n_1160));
   XOR2_X1 i_1201 (.A(n_1160), .B(n_1944), .Z(n_3528));
   INV_X1 i_1202 (.A(n_1117), .ZN(n_1161));
   NAND2_X1 i_1203 (.A1(n_1116), .A2(n_1161), .ZN(n_1162));
   XOR2_X1 i_1204 (.A(n_1162), .B(n_1118), .Z(n_3535));
   INV_X1 i_1205 (.A(n_1126), .ZN(n_1163));
   NAND2_X1 i_1206 (.A1(n_1163), .A2(n_1119), .ZN(n_1166));
   XOR2_X1 i_1207 (.A(n_1166), .B(n_1127), .Z(n_3542));
   INV_X1 i_1210 (.A(n_1132), .ZN(n_1167));
   NAND2_X1 i_1211 (.A1(n_1131), .A2(n_1167), .ZN(n_1168));
   XOR2_X1 i_1212 (.A(n_1168), .B(n_1133), .Z(n_3549));
   INV_X1 i_1213 (.A(n_1136), .ZN(n_1169));
   NAND2_X1 i_1214 (.A1(n_1169), .A2(n_1134), .ZN(n_1170));
   XOR2_X1 i_1215 (.A(n_1170), .B(n_1137), .Z(n_3556));
   INV_X1 i_1216 (.A(n_1140), .ZN(n_1172));
   NAND2_X1 i_1217 (.A1(n_1139), .A2(n_1172), .ZN(n_1173));
   XOR2_X1 i_1218 (.A(n_1173), .B(n_1141), .Z(n_3563));
   INV_X1 i_1219 (.A(n_1145), .ZN(n_1174));
   NAND2_X1 i_1220 (.A1(n_1144), .A2(n_1174), .ZN(n_1175));
   XOR2_X1 i_1221 (.A(n_1175), .B(n_1146), .Z(n_3570));
   NAND4_X1 i_1222 (.A1(in2[21]), .A2(in2[20]), .A3(in1[17]), .A4(in1[16]), 
      .ZN(n_1213));
   AOI22_X1 i_1223 (.A1(in2[21]), .A2(in1[16]), .B1(in2[20]), .B2(in1[17]), 
      .ZN(n_1216));
   NAND2_X1 i_1224 (.A1(in2[22]), .A2(in1[15]), .ZN(n_1217));
   OAI21_X1 i_1225 (.A(n_1213), .B1(n_1216), .B2(n_1217), .ZN(n_3446));
   NAND3_X1 i_1226 (.A1(n_1130), .A2(in1[19]), .A3(in2[18]), .ZN(n_1218));
   AOI21_X1 i_1227 (.A(n_1130), .B1(in1[19]), .B2(in2[18]), .ZN(n_1219));
   NAND2_X1 i_1228 (.A1(in2[19]), .A2(in1[18]), .ZN(n_1220));
   OAI21_X1 i_1229 (.A(n_1218), .B1(n_1219), .B2(n_1220), .ZN(n_3453));
   NAND4_X1 i_1230 (.A1(in1[23]), .A2(in1[22]), .A3(in2[15]), .A4(in2[14]), 
      .ZN(n_1231));
   AOI22_X1 i_1231 (.A1(in1[22]), .A2(in2[15]), .B1(in1[23]), .B2(in2[14]), 
      .ZN(n_1232));
   NAND2_X1 i_1232 (.A1(in1[21]), .A2(in2[16]), .ZN(n_1235));
   OAI21_X1 i_1233 (.A(n_1231), .B1(n_1232), .B2(n_1235), .ZN(n_3460));
   NAND3_X1 i_1234 (.A1(n_1138), .A2(in1[25]), .A3(in2[12]), .ZN(n_1236));
   AOI21_X1 i_1235 (.A(n_1138), .B1(in1[25]), .B2(in2[12]), .ZN(n_1237));
   NAND2_X1 i_1236 (.A1(in1[24]), .A2(in2[13]), .ZN(n_1238));
   OAI21_X1 i_1237 (.A(n_1236), .B1(n_1237), .B2(n_1238), .ZN(n_3467));
   NAND3_X1 i_1238 (.A1(n_1143), .A2(in1[28]), .A3(in2[9]), .ZN(n_1239));
   AOI21_X1 i_1239 (.A(n_1143), .B1(in1[28]), .B2(in2[9]), .ZN(n_1242));
   NAND2_X1 i_1240 (.A1(in1[27]), .A2(in2[10]), .ZN(n_1243));
   OAI21_X1 i_1241 (.A(n_1239), .B1(n_1242), .B2(n_1243), .ZN(n_3474));
   NAND2_X1 i_1242 (.A1(in1[31]), .A2(in2[7]), .ZN(n_516));
   INV_X1 i_1244 (.A(n_1926), .ZN(n_1244));
   NAND2_X1 i_1245 (.A1(n_1244), .A2(n_1927), .ZN(n_1245));
   XOR2_X1 i_1246 (.A(n_1245), .B(n_1925), .Z(n_3422));
   INV_X1 i_1247 (.A(n_1931), .ZN(n_1246));
   NAND2_X1 i_1248 (.A1(n_1932), .A2(n_1246), .ZN(n_1248));
   XOR2_X1 i_1249 (.A(n_1248), .B(n_1930), .Z(n_3431));
   INV_X1 i_1250 (.A(n_1934), .ZN(n_1249));
   NAND2_X1 i_1251 (.A1(n_1937), .A2(n_1249), .ZN(n_1250));
   XOR2_X1 i_1252 (.A(n_1250), .B(n_1933), .Z(n_3438));
   INV_X1 i_1253 (.A(n_1216), .ZN(n_1251));
   NAND2_X1 i_1254 (.A1(n_1251), .A2(n_1213), .ZN(n_1252));
   XOR2_X1 i_1255 (.A(n_1252), .B(n_1217), .Z(n_3445));
   INV_X1 i_1256 (.A(n_1219), .ZN(n_1253));
   NAND2_X1 i_1257 (.A1(n_1218), .A2(n_1253), .ZN(n_1255));
   XOR2_X1 i_1258 (.A(n_1255), .B(n_1220), .Z(n_3452));
   INV_X1 i_1259 (.A(n_1232), .ZN(n_1256));
   NAND2_X1 i_1260 (.A1(n_1256), .A2(n_1231), .ZN(n_1257));
   XOR2_X1 i_1261 (.A(n_1257), .B(n_1235), .Z(n_3459));
   INV_X1 i_1262 (.A(n_1237), .ZN(n_1258));
   NAND2_X1 i_1263 (.A1(n_1236), .A2(n_1258), .ZN(n_1271));
   XOR2_X1 i_1264 (.A(n_1271), .B(n_1238), .Z(n_3466));
   INV_X1 i_1265 (.A(n_1242), .ZN(n_1272));
   NAND2_X1 i_1266 (.A1(n_1239), .A2(n_1272), .ZN(n_1275));
   XOR2_X1 i_1267 (.A(n_1275), .B(n_1243), .Z(n_3473));
   XNOR2_X1 i_1268 (.A(n_1947), .B(n_1953), .ZN(n_3480));
   NAND4_X1 i_1269 (.A1(in2[30]), .A2(in2[29]), .A3(in1[7]), .A4(in1[6]), 
      .ZN(n_1276));
   AOI22_X1 i_1270 (.A1(in2[30]), .A2(in1[6]), .B1(in2[29]), .B2(in1[7]), 
      .ZN(n_1277));
   NOR2_X1 i_1271 (.A1(n_1602), .A2(n_598), .ZN(n_1279));
   OAI21_X1 i_1272 (.A(n_1276), .B1(n_1277), .B2(n_1279), .ZN(n_3324));
   NAND4_X1 i_1273 (.A1(in2[27]), .A2(in2[26]), .A3(in1[10]), .A4(in1[9]), 
      .ZN(n_1282));
   AOI22_X1 i_1274 (.A1(in2[27]), .A2(in1[9]), .B1(in2[26]), .B2(in1[10]), 
      .ZN(n_1283));
   NAND2_X1 i_1275 (.A1(in2[28]), .A2(in1[8]), .ZN(n_1284));
   OAI21_X1 i_1276 (.A(n_1282), .B1(n_1283), .B2(n_1284), .ZN(n_3333));
   INV_X1 i_1277 (.A(n_1277), .ZN(n_1320));
   NAND2_X1 i_1278 (.A1(n_1320), .A2(n_1276), .ZN(n_1323));
   XOR2_X1 i_1279 (.A(n_1323), .B(n_1279), .Z(n_3323));
   INV_X1 i_1280 (.A(n_1283), .ZN(n_1324));
   NAND2_X1 i_1281 (.A1(n_1324), .A2(n_1282), .ZN(n_1325));
   XOR2_X1 i_1282 (.A(n_1325), .B(n_1284), .Z(n_3332));
   INV_X1 i_1283 (.A(n_2000), .ZN(n_1326));
   NAND2_X1 i_1284 (.A1(n_1326), .A2(n_2001), .ZN(n_1327));
   XOR2_X1 i_1286 (.A(n_1327), .B(n_1999), .Z(n_3339));
   INV_X1 i_1287 (.A(n_2003), .ZN(n_1330));
   NAND2_X1 i_1288 (.A1(n_1330), .A2(n_2070), .ZN(n_1331));
   XOR2_X1 i_1289 (.A(n_1331), .B(n_2002), .Z(n_3346));
   INV_X1 i_1290 (.A(n_2072), .ZN(n_1332));
   NAND2_X1 i_1291 (.A1(n_1332), .A2(n_2073), .ZN(n_1333));
   XOR2_X1 i_1292 (.A(n_1333), .B(n_2071), .Z(n_3353));
   INV_X1 i_1293 (.A(n_1987), .ZN(n_1334));
   NAND2_X1 i_1294 (.A1(n_1334), .A2(n_1988), .ZN(n_1337));
   XOR2_X1 i_1295 (.A(n_1337), .B(n_1986), .Z(n_3360));
   INV_X1 i_1296 (.A(n_1992), .ZN(n_1338));
   NAND2_X1 i_1297 (.A1(n_1338), .A2(n_1993), .ZN(n_1339));
   XOR2_X1 i_1298 (.A(n_1339), .B(n_1989), .Z(n_3367));
   INV_X1 i_1299 (.A(n_1995), .ZN(n_1340));
   NAND2_X1 i_1300 (.A1(n_1340), .A2(n_1996), .ZN(n_1341));
   XOR2_X1 i_1301 (.A(n_1341), .B(n_1994), .Z(n_3374));
   NAND2_X1 i_1302 (.A1(n_1985), .A2(n_1982), .ZN(n_1344));
   XOR2_X1 i_1303 (.A(n_1344), .B(n_1954), .Z(n_3380));
   NAND4_X1 i_1304 (.A1(in1[23]), .A2(in1[24]), .A3(in2[12]), .A4(in2[11]), 
      .ZN(n_1388));
   AOI22_X1 i_1305 (.A1(in1[23]), .A2(in2[12]), .B1(in1[24]), .B2(in2[11]), 
      .ZN(n_1389));
   NAND2_X1 i_1306 (.A1(in1[22]), .A2(in2[13]), .ZN(n_1390));
   OAI21_X1 i_1307 (.A(n_1388), .B1(n_1389), .B2(n_1390), .ZN(n_3268));
   NAND4_X1 i_1308 (.A1(in1[26]), .A2(in1[27]), .A3(in2[9]), .A4(in2[8]), 
      .ZN(n_1391));
   AOI22_X1 i_1309 (.A1(in1[26]), .A2(in2[9]), .B1(in1[27]), .B2(in2[8]), 
      .ZN(n_1393));
   NAND2_X1 i_1310 (.A1(in1[25]), .A2(in2[10]), .ZN(n_1394));
   OAI21_X1 i_1311 (.A(n_1391), .B1(n_1393), .B2(n_1394), .ZN(n_3275));
   NAND4_X1 i_1312 (.A1(in1[29]), .A2(in1[30]), .A3(in2[6]), .A4(in2[5]), 
      .ZN(n_1395));
   AOI22_X1 i_1313 (.A1(in1[29]), .A2(in2[6]), .B1(in1[30]), .B2(in2[5]), 
      .ZN(n_1396));
   NAND2_X1 i_1314 (.A1(in1[28]), .A2(in2[7]), .ZN(n_1397));
   OAI21_X1 i_1315 (.A(n_1395), .B1(n_1396), .B2(n_1397), .ZN(n_3282));
   INV_X1 i_1316 (.A(n_1856), .ZN(n_1398));
   NAND2_X1 i_1317 (.A1(n_1853), .A2(n_1398), .ZN(n_1400));
   XOR2_X1 i_1318 (.A(n_1400), .B(n_1858), .Z(n_3223));
   INV_X1 i_1319 (.A(n_1860), .ZN(n_1401));
   NAND2_X1 i_1320 (.A1(n_1401), .A2(n_1859), .ZN(n_1402));
   XOR2_X1 i_1321 (.A(n_1402), .B(n_1862), .Z(n_3232));
   INV_X1 i_1322 (.A(n_1864), .ZN(n_1403));
   NAND2_X1 i_1323 (.A1(n_1403), .A2(n_1863), .ZN(n_1420));
   XOR2_X1 i_1324 (.A(n_1420), .B(n_1865), .Z(n_3239));
   INV_X1 i_1325 (.A(n_1843), .ZN(n_1421));
   NAND2_X1 i_1326 (.A1(n_1421), .A2(n_1842), .ZN(n_1424));
   XOR2_X1 i_1327 (.A(n_1424), .B(n_1844), .Z(n_3246));
   INV_X1 i_1328 (.A(n_1846), .ZN(n_1425));
   NAND2_X1 i_1329 (.A1(n_1425), .A2(n_1845), .ZN(n_1426));
   XOR2_X1 i_1330 (.A(n_1426), .B(n_1849), .Z(n_3253));
   INV_X1 i_1331 (.A(n_1851), .ZN(n_1427));
   NAND2_X1 i_1332 (.A1(n_1427), .A2(n_1850), .ZN(n_1428));
   XOR2_X1 i_1333 (.A(n_1428), .B(n_1852), .Z(n_3260));
   INV_X1 i_1334 (.A(n_1389), .ZN(n_1431));
   NAND2_X1 i_1335 (.A1(n_1431), .A2(n_1388), .ZN(n_1432));
   XOR2_X1 i_1336 (.A(n_1432), .B(n_1390), .Z(n_3267));
   INV_X1 i_1337 (.A(n_1393), .ZN(n_1433));
   NAND2_X1 i_1338 (.A1(n_1433), .A2(n_1391), .ZN(n_1434));
   XOR2_X1 i_1339 (.A(n_1434), .B(n_1394), .Z(n_3274));
   INV_X1 i_1340 (.A(n_1396), .ZN(n_1435));
   NAND2_X1 i_1341 (.A1(n_1435), .A2(n_1395), .ZN(n_1438));
   XOR2_X1 i_1342 (.A(n_1438), .B(n_1397), .Z(n_3281));
   OAI21_X1 i_1343 (.A(n_1683), .B1(n_1678), .B2(n_1679), .ZN(n_1453));
   INV_X1 i_1344 (.A(n_1678), .ZN(n_1454));
   OAI21_X1 i_1345 (.A(n_1453), .B1(n_1454), .B2(n_1680), .ZN(n_3181));
   NAND2_X1 i_1346 (.A1(n_1872), .A2(n_1904), .ZN(n_1552));
   XOR2_X1 i_1347 (.A(n_1552), .B(n_1905), .Z(n_3115));
   NOR2_X1 i_1348 (.A1(n_1831), .A2(n_1830), .ZN(n_1783));
   XNOR2_X1 i_1349 (.A(n_1783), .B(n_1375), .ZN(n_2932));
   NOR2_X1 i_1350 (.A1(n_1791), .A2(n_1782), .ZN(n_1784));
   XNOR2_X1 i_1351 (.A(n_1784), .B(n_1305), .ZN(n_2939));
   NOR2_X1 i_1352 (.A1(n_1825), .A2(n_1824), .ZN(n_1785));
   XNOR2_X1 i_1353 (.A(n_1785), .B(n_1345), .ZN(n_2946));
   NOR2_X1 i_1354 (.A1(n_1829), .A2(n_1828), .ZN(n_1786));
   XNOR2_X1 i_1355 (.A(n_1786), .B(n_1350), .ZN(n_2953));
   NAND2_X1 i_1356 (.A1(n_1286), .A2(n_1204), .ZN(n_1787));
   XOR2_X1 i_1357 (.A(n_1205), .B(n_1787), .Z(n_2960));
   OAI211_X1 i_1358 (.A(in1[31]), .B(in2[0]), .C1(n_1383), .C2(n_1377), .ZN(
      n_1789));
   INV_X1 i_1359 (.A(n_1789), .ZN(n_1790));
   NAND3_X1 i_1360 (.A1(n_1514), .A2(in1[29]), .A3(in2[2]), .ZN(n_1792));
   INV_X1 i_1361 (.A(n_1792), .ZN(n_1817));
   NOR2_X1 i_1362 (.A1(n_1381), .A2(n_599), .ZN(n_1818));
   OAI21_X1 i_1363 (.A(n_1278), .B1(n_1382), .B2(n_1377), .ZN(n_1821));
   AOI21_X1 i_1364 (.A(n_1817), .B1(n_1818), .B2(n_1821), .ZN(n_1822));
   OAI211_X1 i_1365 (.A(in1[30]), .B(in2[1]), .C1(n_1384), .C2(n_692), .ZN(
      n_1823));
   AOI21_X1 i_1366 (.A(n_1790), .B1(n_1822), .B2(n_1823), .ZN(n_2848));
   INV_X1 i_1367 (.A(n_1566), .ZN(n_1873));
   NAND2_X1 i_1368 (.A1(n_1567), .A2(n_1873), .ZN(n_1898));
   XOR2_X1 i_1369 (.A(n_1898), .B(n_1565), .Z(n_2775));
   INV_X1 i_1370 (.A(n_1571), .ZN(n_1899));
   NAND2_X1 i_1371 (.A1(n_1572), .A2(n_1899), .ZN(n_1902));
   XOR2_X1 i_1372 (.A(n_1902), .B(n_1569), .Z(n_2784));
   INV_X1 i_1373 (.A(n_1299), .ZN(n_1919));
   NAND2_X1 i_1374 (.A1(n_1300), .A2(n_1919), .ZN(n_1920));
   XOR2_X1 i_1375 (.A(n_1920), .B(n_1298), .Z(n_2833));
   NAND2_X1 i_1376 (.A1(n_1211), .A2(n_1206), .ZN(n_1923));
   XNOR2_X1 i_1377 (.A(n_1923), .B(n_1210), .ZN(n_2840));
   NAND2_X1 i_1378 (.A1(n_1789), .A2(n_1823), .ZN(n_1924));
   XOR2_X1 i_1379 (.A(n_1822), .B(n_1924), .Z(n_2847));
   INV_X1 i_1380 (.A(n_1501), .ZN(n_2006));
   NAND2_X1 i_1381 (.A1(n_1499), .A2(n_2006), .ZN(n_2007));
   XOR2_X1 i_1382 (.A(n_2007), .B(n_1500), .Z(n_2732));
   INV_X1 i_1383 (.A(n_1771), .ZN(n_2008));
   NAND2_X1 i_1384 (.A1(n_1772), .A2(n_2008), .ZN(n_2009));
   XOR2_X1 i_1385 (.A(n_2009), .B(n_1770), .Z(n_2662));
   INV_X1 i_1386 (.A(n_1776), .ZN(n_2010));
   NAND2_X1 i_1387 (.A1(n_1777), .A2(n_2010), .ZN(n_2013));
   XOR2_X1 i_1388 (.A(n_2013), .B(n_1773), .Z(n_2669));
   INV_X1 i_1389 (.A(n_1779), .ZN(n_2014));
   NAND2_X1 i_1390 (.A1(n_2014), .A2(n_1780), .ZN(n_2015));
   XOR2_X1 i_1391 (.A(n_2015), .B(n_1778), .Z(n_2676));
   INV_X1 i_1392 (.A(n_1758), .ZN(n_2016));
   NAND2_X1 i_1393 (.A1(n_2016), .A2(n_1759), .ZN(n_2017));
   XOR2_X1 i_1394 (.A(n_2017), .B(n_1757), .Z(n_2683));
   INV_X1 i_1395 (.A(n_1763), .ZN(n_2020));
   NAND2_X1 i_1396 (.A1(n_2020), .A2(n_1764), .ZN(n_2021));
   XOR2_X1 i_1397 (.A(n_2021), .B(n_1762), .Z(n_2690));
   INV_X1 i_1398 (.A(n_1766), .ZN(n_2022));
   NAND2_X1 i_1399 (.A1(n_2022), .A2(n_1769), .ZN(n_2023));
   XOR2_X1 i_1400 (.A(n_2023), .B(n_1765), .Z(n_2697));
   INV_X1 i_1401 (.A(n_1745), .ZN(n_2024));
   NAND2_X1 i_1402 (.A1(n_2024), .A2(n_1748), .ZN(n_2026));
   XOR2_X1 i_1403 (.A(n_2026), .B(n_1744), .Z(n_2704));
   INV_X1 i_1404 (.A(n_1750), .ZN(n_2027));
   NAND2_X1 i_1405 (.A1(n_2027), .A2(n_1751), .ZN(n_2028));
   XOR2_X1 i_1406 (.A(n_2028), .B(n_1749), .Z(n_2711));
   INV_X1 i_1407 (.A(n_1755), .ZN(n_2029));
   NAND2_X1 i_1408 (.A1(n_2029), .A2(n_1756), .ZN(n_2030));
   XOR2_X1 i_1409 (.A(n_2030), .B(n_1752), .Z(n_2718));
   NAND2_X1 i_1410 (.A1(n_1792), .A2(n_1821), .ZN(n_2031));
   XNOR2_X1 i_1411 (.A(n_2031), .B(n_1818), .ZN(n_2725));
   NAND4_X1 i_1412 (.A1(in2[28]), .A2(in2[27]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2033));
   AOI22_X1 i_1413 (.A1(in2[27]), .A2(in1[2]), .B1(in2[28]), .B2(in1[1]), 
      .ZN(n_2034));
   NAND2_X1 i_1414 (.A1(in2[29]), .A2(in1[0]), .ZN(n_2035));
   OAI21_X1 i_1415 (.A(n_2033), .B1(n_2034), .B2(n_2035), .ZN(n_2557));
   NOR2_X1 i_1416 (.A1(n_3574), .A2(n_598), .ZN(n_2036));
   NAND3_X1 i_1417 (.A1(n_2036), .A2(in2[25]), .A3(in1[4]), .ZN(n_2065));
   AOI21_X1 i_1418 (.A(n_2036), .B1(in2[25]), .B2(in1[4]), .ZN(n_2066));
   NAND2_X1 i_1419 (.A1(in2[26]), .A2(in1[3]), .ZN(n_2069));
   OAI21_X1 i_1420 (.A(n_2065), .B1(n_2066), .B2(n_2069), .ZN(n_2564));
   INV_X1 i_1421 (.A(n_2034), .ZN(n_2094));
   NAND2_X1 i_1422 (.A1(n_2094), .A2(n_2033), .ZN(n_2097));
   XOR2_X1 i_1423 (.A(n_2097), .B(n_2035), .Z(n_2556));
   INV_X1 i_1424 (.A(n_2066), .ZN(n_2098));
   NAND2_X1 i_1425 (.A1(n_2065), .A2(n_2098), .ZN(n_2099));
   XOR2_X1 i_1426 (.A(n_2099), .B(n_2069), .Z(n_2563));
   INV_X1 i_1427 (.A(n_1547), .ZN(n_2100));
   NAND2_X1 i_1428 (.A1(n_2100), .A2(n_1548), .ZN(n_2101));
   XOR2_X1 i_1429 (.A(n_2101), .B(n_1546), .Z(n_2570));
   INV_X1 i_1430 (.A(n_1553), .ZN(n_2104));
   NAND2_X1 i_1431 (.A1(n_2104), .A2(n_1554), .ZN(n_2105));
   XOR2_X1 i_1432 (.A(n_2105), .B(n_1551), .Z(n_2577));
   INV_X1 i_1433 (.A(n_1558), .ZN(n_2106));
   NAND2_X1 i_1434 (.A1(n_2106), .A2(n_1559), .ZN(n_2107));
   XOR2_X1 i_1435 (.A(n_2107), .B(n_1555), .Z(n_2584));
   INV_X1 i_1436 (.A(n_1518), .ZN(n_2108));
   NAND2_X1 i_1437 (.A1(n_2108), .A2(n_1519), .ZN(n_2111));
   XOR2_X1 i_1438 (.A(n_2111), .B(n_1517), .Z(n_2591));
   INV_X1 i_1439 (.A(n_1521), .ZN(n_2112));
   NAND2_X1 i_1440 (.A1(n_2112), .A2(n_1540), .ZN(n_2113));
   XOR2_X1 i_1441 (.A(n_2113), .B(n_1520), .Z(n_2598));
   INV_X1 i_1442 (.A(n_1544), .ZN(n_2114));
   NAND2_X1 i_1443 (.A1(n_2114), .A2(n_1545), .ZN(n_2115));
   XOR2_X1 i_1444 (.A(n_2115), .B(n_1541), .Z(n_2605));
   INV_X1 i_1445 (.A(n_1507), .ZN(n_2117));
   NAND2_X1 i_1446 (.A1(n_2117), .A2(n_1508), .ZN(n_2118));
   XOR2_X1 i_1447 (.A(n_2118), .B(n_1506), .Z(n_2612));
   INV_X1 i_1448 (.A(n_1512), .ZN(n_2119));
   NAND2_X1 i_1449 (.A1(n_1513), .A2(n_2119), .ZN(n_2120));
   XOR2_X1 i_1450 (.A(n_2120), .B(n_1511), .Z(n_2619));
   NAND4_X1 i_1451 (.A1(in1[26]), .A2(in1[25]), .A3(in2[2]), .A4(in2[1]), 
      .ZN(n_2121));
   AOI22_X1 i_1452 (.A1(in1[26]), .A2(in2[1]), .B1(in1[25]), .B2(in2[2]), 
      .ZN(n_2122));
   NAND2_X1 i_1453 (.A1(in1[24]), .A2(in2[3]), .ZN(n_2125));
   OAI21_X1 i_1454 (.A(n_2121), .B1(n_2122), .B2(n_2125), .ZN(n_2126));
   AOI21_X1 i_1455 (.A(n_2126), .B1(in1[28]), .B2(in2[0]), .ZN(n_2127));
   NAND2_X1 i_1456 (.A1(in1[27]), .A2(in2[1]), .ZN(n_2128));
   NAND3_X1 i_1457 (.A1(n_2126), .A2(in1[28]), .A3(in2[0]), .ZN(n_2157));
   AOI21_X1 i_1458 (.A(n_2127), .B1(n_2128), .B2(n_2157), .ZN(n_2514));
   NAND4_X1 i_1459 (.A1(in2[27]), .A2(in2[26]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2158));
   AOI22_X1 i_1460 (.A1(in2[26]), .A2(in1[2]), .B1(in2[27]), .B2(in1[1]), 
      .ZN(n_2161));
   NAND2_X1 i_1461 (.A1(in2[28]), .A2(in1[0]), .ZN(n_2162));
   OAI21_X1 i_1462 (.A(n_2158), .B1(n_2161), .B2(n_2162), .ZN(n_2452));
   NOR2_X1 i_1463 (.A1(n_3649), .A2(n_598), .ZN(n_2163));
   NAND3_X1 i_1464 (.A1(n_2163), .A2(in2[24]), .A3(in1[4]), .ZN(n_2164));
   AOI21_X1 i_1465 (.A(n_2163), .B1(in2[24]), .B2(in1[4]), .ZN(n_2165));
   NAND2_X1 i_1466 (.A1(in2[25]), .A2(in1[3]), .ZN(n_2168));
   OAI21_X1 i_1467 (.A(n_2164), .B1(n_2165), .B2(n_2168), .ZN(n_2459));
   NAND4_X1 i_1468 (.A1(in2[21]), .A2(in2[20]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2169));
   AOI22_X1 i_1469 (.A1(in2[20]), .A2(in1[8]), .B1(in2[21]), .B2(in1[7]), 
      .ZN(n_2170));
   NAND2_X1 i_1470 (.A1(in2[22]), .A2(in1[6]), .ZN(n_2171));
   OAI21_X1 i_1471 (.A(n_2169), .B1(n_2170), .B2(n_2171), .ZN(n_2466));
   NAND4_X1 i_1472 (.A1(in2[18]), .A2(in2[17]), .A3(in1[11]), .A4(in1[10]), 
      .ZN(n_2172));
   AOI22_X1 i_1473 (.A1(in2[17]), .A2(in1[11]), .B1(in2[18]), .B2(in1[10]), 
      .ZN(n_2175));
   NAND2_X1 i_1474 (.A1(in2[19]), .A2(in1[9]), .ZN(n_2176));
   OAI21_X1 i_1475 (.A(n_2172), .B1(n_2175), .B2(n_2176), .ZN(n_2473));
   NAND4_X1 i_1476 (.A1(in1[14]), .A2(in2[15]), .A3(in2[14]), .A4(in1[13]), 
      .ZN(n_2177));
   AOI22_X1 i_1477 (.A1(in1[14]), .A2(in2[14]), .B1(in2[15]), .B2(in1[13]), 
      .ZN(n_2178));
   NAND2_X1 i_1478 (.A1(in2[16]), .A2(in1[12]), .ZN(n_2179));
   OAI21_X1 i_1479 (.A(n_2177), .B1(n_2178), .B2(n_2179), .ZN(n_2480));
   NAND4_X1 i_1480 (.A1(in1[17]), .A2(in1[16]), .A3(in2[12]), .A4(in2[11]), 
      .ZN(n_2182));
   AOI22_X1 i_1481 (.A1(in1[17]), .A2(in2[11]), .B1(in1[16]), .B2(in2[12]), 
      .ZN(n_2183));
   NAND2_X1 i_1482 (.A1(in1[15]), .A2(in2[13]), .ZN(n_2184));
   OAI21_X1 i_1483 (.A(n_2182), .B1(n_2183), .B2(n_2184), .ZN(n_2487));
   NAND4_X1 i_1484 (.A1(in1[20]), .A2(in1[19]), .A3(in2[9]), .A4(in2[8]), 
      .ZN(n_2185));
   AOI22_X1 i_1485 (.A1(in1[20]), .A2(in2[8]), .B1(in1[19]), .B2(in2[9]), 
      .ZN(n_2186));
   NAND2_X1 i_1486 (.A1(in1[18]), .A2(in2[10]), .ZN(n_2189));
   OAI21_X1 i_1487 (.A(n_2185), .B1(n_2186), .B2(n_2189), .ZN(n_2494));
   NAND4_X1 i_1488 (.A1(in1[23]), .A2(in1[22]), .A3(in2[6]), .A4(in2[5]), 
      .ZN(n_2190));
   AOI22_X1 i_1489 (.A1(in1[23]), .A2(in2[5]), .B1(in1[22]), .B2(in2[6]), 
      .ZN(n_2191));
   NAND2_X1 i_1490 (.A1(in1[21]), .A2(in2[7]), .ZN(n_2192));
   OAI21_X1 i_1491 (.A(n_2190), .B1(n_2191), .B2(n_2192), .ZN(n_2501));
   NAND4_X1 i_1492 (.A1(in1[26]), .A2(in1[25]), .A3(in2[2]), .A4(in2[3]), 
      .ZN(n_2193));
   AOI22_X1 i_1493 (.A1(in1[26]), .A2(in2[2]), .B1(in1[25]), .B2(in2[3]), 
      .ZN(n_2196));
   NAND2_X1 i_1494 (.A1(in1[24]), .A2(in2[4]), .ZN(n_2197));
   OAI21_X1 i_1495 (.A(n_2193), .B1(n_2196), .B2(n_2197), .ZN(n_2508));
   INV_X1 i_1496 (.A(n_2161), .ZN(n_2198));
   NAND2_X1 i_1497 (.A1(n_2198), .A2(n_2158), .ZN(n_2199));
   XOR2_X1 i_1498 (.A(n_2199), .B(n_2162), .Z(n_2451));
   INV_X1 i_1499 (.A(n_2165), .ZN(n_2200));
   NAND2_X1 i_1500 (.A1(n_2164), .A2(n_2200), .ZN(n_2203));
   XOR2_X1 i_1501 (.A(n_2203), .B(n_2168), .Z(n_2458));
   INV_X1 i_1502 (.A(n_2170), .ZN(n_2204));
   NAND2_X1 i_1503 (.A1(n_2204), .A2(n_2169), .ZN(n_2205));
   XOR2_X1 i_1504 (.A(n_2205), .B(n_2171), .Z(n_2465));
   INV_X1 i_1505 (.A(n_2175), .ZN(n_2206));
   NAND2_X1 i_1506 (.A1(n_2206), .A2(n_2172), .ZN(n_2207));
   XOR2_X1 i_1507 (.A(n_2207), .B(n_2176), .Z(n_2472));
   INV_X1 i_1508 (.A(n_2178), .ZN(n_2210));
   NAND2_X1 i_1509 (.A1(n_2210), .A2(n_2177), .ZN(n_2211));
   XOR2_X1 i_1510 (.A(n_2211), .B(n_2179), .Z(n_2479));
   INV_X1 i_1511 (.A(n_2183), .ZN(n_2212));
   NAND2_X1 i_1512 (.A1(n_2212), .A2(n_2182), .ZN(n_2213));
   XOR2_X1 i_1513 (.A(n_2213), .B(n_2184), .Z(n_2486));
   INV_X1 i_1514 (.A(n_2186), .ZN(n_2216));
   NAND2_X1 i_1515 (.A1(n_2216), .A2(n_2185), .ZN(n_2217));
   XOR2_X1 i_1516 (.A(n_2217), .B(n_2189), .Z(n_2493));
   INV_X1 i_1517 (.A(n_2191), .ZN(n_2218));
   NAND2_X1 i_1518 (.A1(n_2218), .A2(n_2190), .ZN(n_2219));
   XOR2_X1 i_1519 (.A(n_2219), .B(n_2192), .Z(n_2500));
   INV_X1 i_1520 (.A(n_2196), .ZN(n_2220));
   NAND2_X1 i_1521 (.A1(n_2220), .A2(n_2193), .ZN(n_2251));
   XOR2_X1 i_1522 (.A(n_2251), .B(n_2197), .Z(n_2507));
   INV_X1 i_1523 (.A(n_2127), .ZN(n_2252));
   NAND2_X1 i_1524 (.A1(n_2252), .A2(n_2157), .ZN(n_2255));
   XOR2_X1 i_1525 (.A(n_2255), .B(n_2128), .Z(n_2513));
   NAND2_X1 i_1526 (.A1(in1[27]), .A2(in2[0]), .ZN(n_2269));
   AOI21_X1 i_1527 (.A(n_697), .B1(n_2269), .B2(n_696), .ZN(n_2412));
   NAND4_X1 i_1528 (.A1(in2[26]), .A2(in2[25]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2271));
   AOI22_X1 i_1529 (.A1(in2[25]), .A2(in1[2]), .B1(in2[26]), .B2(in1[1]), 
      .ZN(n_2272));
   NAND2_X1 i_1530 (.A1(in2[27]), .A2(in1[0]), .ZN(n_2273));
   OAI21_X1 i_1531 (.A(n_2271), .B1(n_2272), .B2(n_2273), .ZN(n_2349));
   NAND3_X1 i_1532 (.A1(n_2163), .A2(in2[22]), .A3(in1[4]), .ZN(n_2276));
   AOI22_X1 i_1533 (.A1(in2[22]), .A2(in1[5]), .B1(in2[23]), .B2(in1[4]), 
      .ZN(n_2277));
   NAND2_X1 i_1534 (.A1(in2[24]), .A2(in1[3]), .ZN(n_2278));
   OAI21_X1 i_1535 (.A(n_2276), .B1(n_2277), .B2(n_2278), .ZN(n_2356));
   NAND4_X1 i_1536 (.A1(in2[20]), .A2(in2[19]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2279));
   AOI22_X1 i_1537 (.A1(in2[19]), .A2(in1[8]), .B1(in2[20]), .B2(in1[7]), 
      .ZN(n_2280));
   NAND2_X1 i_1538 (.A1(in2[21]), .A2(in1[6]), .ZN(n_2283));
   OAI21_X1 i_1539 (.A(n_2279), .B1(n_2280), .B2(n_2283), .ZN(n_2363));
   NAND4_X1 i_1540 (.A1(in2[17]), .A2(in2[16]), .A3(in1[11]), .A4(in1[10]), 
      .ZN(n_2284));
   AOI22_X1 i_1541 (.A1(in2[16]), .A2(in1[11]), .B1(in2[17]), .B2(in1[10]), 
      .ZN(n_2285));
   NAND2_X1 i_1542 (.A1(in2[18]), .A2(in1[9]), .ZN(n_2286));
   OAI21_X1 i_1543 (.A(n_2284), .B1(n_2285), .B2(n_2286), .ZN(n_2370));
   NAND4_X1 i_1544 (.A1(in1[14]), .A2(in2[14]), .A3(in1[13]), .A4(in2[13]), 
      .ZN(n_2287));
   AOI22_X1 i_1545 (.A1(in1[14]), .A2(in2[13]), .B1(in2[14]), .B2(in1[13]), 
      .ZN(n_2290));
   NAND2_X1 i_1546 (.A1(in2[15]), .A2(in1[12]), .ZN(n_2291));
   OAI21_X1 i_1547 (.A(n_2287), .B1(n_2290), .B2(n_2291), .ZN(n_2377));
   NAND4_X1 i_1548 (.A1(in1[17]), .A2(in1[16]), .A3(in2[11]), .A4(in2[10]), 
      .ZN(n_2292));
   AOI22_X1 i_1549 (.A1(in1[17]), .A2(in2[10]), .B1(in1[16]), .B2(in2[11]), 
      .ZN(n_2293));
   NAND2_X1 i_1550 (.A1(in1[15]), .A2(in2[12]), .ZN(n_2294));
   OAI21_X1 i_1551 (.A(n_2292), .B1(n_2293), .B2(n_2294), .ZN(n_2384));
   NAND4_X1 i_1552 (.A1(in1[20]), .A2(in1[19]), .A3(in2[8]), .A4(in2[7]), 
      .ZN(n_2297));
   AOI22_X1 i_1553 (.A1(in1[20]), .A2(in2[7]), .B1(in1[19]), .B2(in2[8]), 
      .ZN(n_2298));
   NAND2_X1 i_1554 (.A1(in1[18]), .A2(in2[9]), .ZN(n_2299));
   OAI21_X1 i_1555 (.A(n_2297), .B1(n_2298), .B2(n_2299), .ZN(n_2391));
   NAND4_X1 i_1556 (.A1(in1[23]), .A2(in1[22]), .A3(in2[4]), .A4(in2[5]), 
      .ZN(n_2300));
   AOI22_X1 i_1557 (.A1(in1[23]), .A2(in2[4]), .B1(in1[22]), .B2(in2[5]), 
      .ZN(n_2301));
   NAND2_X1 i_1558 (.A1(in1[21]), .A2(in2[6]), .ZN(n_2303));
   OAI21_X1 i_1559 (.A(n_2300), .B1(n_2301), .B2(n_2303), .ZN(n_2398));
   XOR2_X1 i_1560 (.A(n_695), .B(n_2269), .Z(n_2411));
   INV_X1 i_1561 (.A(n_2272), .ZN(n_2306));
   NAND2_X1 i_1562 (.A1(n_2306), .A2(n_2271), .ZN(n_2307));
   XOR2_X1 i_1563 (.A(n_2307), .B(n_2273), .Z(n_2348));
   INV_X1 i_1564 (.A(n_2277), .ZN(n_2308));
   NAND2_X1 i_1565 (.A1(n_2276), .A2(n_2308), .ZN(n_2310));
   XOR2_X1 i_1566 (.A(n_2310), .B(n_2278), .Z(n_2355));
   INV_X1 i_1567 (.A(n_2280), .ZN(n_2311));
   NAND2_X1 i_1568 (.A1(n_2311), .A2(n_2279), .ZN(n_2312));
   XOR2_X1 i_1569 (.A(n_2312), .B(n_2283), .Z(n_2362));
   INV_X1 i_1570 (.A(n_2285), .ZN(n_2313));
   NAND2_X1 i_1571 (.A1(n_2313), .A2(n_2284), .ZN(n_2346));
   XOR2_X1 i_1572 (.A(n_2346), .B(n_2286), .Z(n_2369));
   INV_X1 i_1573 (.A(n_2290), .ZN(n_2347));
   NAND2_X1 i_1574 (.A1(n_2347), .A2(n_2287), .ZN(n_2350));
   XOR2_X1 i_1575 (.A(n_2350), .B(n_2291), .Z(n_2376));
   INV_X1 i_1576 (.A(n_2293), .ZN(n_2351));
   NAND2_X1 i_1577 (.A1(n_2351), .A2(n_2292), .ZN(n_2352));
   XOR2_X1 i_1578 (.A(n_2352), .B(n_2294), .Z(n_2383));
   INV_X1 i_1579 (.A(n_2298), .ZN(n_2353));
   NAND2_X1 i_1580 (.A1(n_2353), .A2(n_2297), .ZN(n_2354));
   XOR2_X1 i_1581 (.A(n_2354), .B(n_2299), .Z(n_2390));
   INV_X1 i_1582 (.A(n_2301), .ZN(n_2357));
   NAND2_X1 i_1583 (.A1(n_2357), .A2(n_2300), .ZN(n_2358));
   XOR2_X1 i_1584 (.A(n_2358), .B(n_2303), .Z(n_2397));
   INV_X1 i_1585 (.A(n_2122), .ZN(n_2359));
   NAND2_X1 i_1586 (.A1(n_2359), .A2(n_2121), .ZN(n_2360));
   XOR2_X1 i_1587 (.A(n_2360), .B(n_2125), .Z(n_2404));
   NAND4_X1 i_1588 (.A1(in2[25]), .A2(in2[24]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2361));
   AOI22_X1 i_1589 (.A1(in2[24]), .A2(in1[2]), .B1(in2[25]), .B2(in1[1]), 
      .ZN(n_2364));
   NAND2_X1 i_1590 (.A1(in2[26]), .A2(in1[0]), .ZN(n_2365));
   OAI21_X1 i_1591 (.A(n_2361), .B1(n_2364), .B2(n_2365), .ZN(n_2254));
   NOR2_X1 i_1592 (.A1(n_3573), .A2(n_598), .ZN(n_2366));
   NAND3_X1 i_1593 (.A1(n_2366), .A2(in2[22]), .A3(in1[4]), .ZN(n_2367));
   AOI21_X1 i_1594 (.A(n_2366), .B1(in2[22]), .B2(in1[4]), .ZN(n_2368));
   NAND2_X1 i_1595 (.A1(in2[23]), .A2(in1[3]), .ZN(n_2371));
   OAI21_X1 i_1596 (.A(n_2367), .B1(n_2368), .B2(n_2371), .ZN(n_2261));
   NAND4_X1 i_1597 (.A1(in2[19]), .A2(in2[18]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2372));
   AOI22_X1 i_1598 (.A1(in2[18]), .A2(in1[8]), .B1(in2[19]), .B2(in1[7]), 
      .ZN(n_2373));
   NAND2_X1 i_1599 (.A1(in2[20]), .A2(in1[6]), .ZN(n_2374));
   OAI21_X1 i_1600 (.A(n_2372), .B1(n_2373), .B2(n_2374), .ZN(n_2268));
   NAND4_X1 i_1601 (.A1(in2[16]), .A2(in2[15]), .A3(in1[11]), .A4(in1[10]), 
      .ZN(n_2375));
   AOI22_X1 i_1602 (.A1(in2[15]), .A2(in1[11]), .B1(in2[16]), .B2(in1[10]), 
      .ZN(n_2378));
   NAND2_X1 i_1603 (.A1(in2[17]), .A2(in1[9]), .ZN(n_2379));
   OAI21_X1 i_1604 (.A(n_2375), .B1(n_2378), .B2(n_2379), .ZN(n_2275));
   NAND4_X1 i_1605 (.A1(in1[14]), .A2(in1[13]), .A3(in2[13]), .A4(in2[12]), 
      .ZN(n_2380));
   AOI22_X1 i_1606 (.A1(in1[14]), .A2(in2[12]), .B1(in1[13]), .B2(in2[13]), 
      .ZN(n_2381));
   NAND2_X1 i_1607 (.A1(in2[14]), .A2(in1[12]), .ZN(n_2382));
   OAI21_X1 i_1608 (.A(n_2380), .B1(n_2381), .B2(n_2382), .ZN(n_2282));
   NAND4_X1 i_1609 (.A1(in1[17]), .A2(in1[16]), .A3(in2[10]), .A4(in2[9]), 
      .ZN(n_2385));
   AOI22_X1 i_1610 (.A1(in1[17]), .A2(in2[9]), .B1(in1[16]), .B2(in2[10]), 
      .ZN(n_2386));
   NAND2_X1 i_1611 (.A1(in1[15]), .A2(in2[11]), .ZN(n_2387));
   OAI21_X1 i_1612 (.A(n_2385), .B1(n_2386), .B2(n_2387), .ZN(n_2289));
   NAND4_X1 i_1613 (.A1(in1[20]), .A2(in1[19]), .A3(in2[7]), .A4(in2[6]), 
      .ZN(n_2388));
   AOI22_X1 i_1614 (.A1(in1[20]), .A2(in2[6]), .B1(in1[19]), .B2(in2[7]), 
      .ZN(n_2389));
   NAND2_X1 i_1615 (.A1(in1[18]), .A2(in2[8]), .ZN(n_2392));
   OAI21_X1 i_1616 (.A(n_2388), .B1(n_2389), .B2(n_2392), .ZN(n_2296));
   INV_X1 i_1617 (.A(n_2364), .ZN(n_2393));
   NAND2_X1 i_1618 (.A1(n_2393), .A2(n_2361), .ZN(n_2394));
   XOR2_X1 i_1619 (.A(n_2394), .B(n_2365), .Z(n_2253));
   INV_X1 i_1620 (.A(n_2368), .ZN(n_2395));
   NAND2_X1 i_1621 (.A1(n_2367), .A2(n_2395), .ZN(n_2396));
   XOR2_X1 i_1622 (.A(n_2396), .B(n_2371), .Z(n_2260));
   INV_X1 i_1623 (.A(n_2373), .ZN(n_2399));
   NAND2_X1 i_1624 (.A1(n_2399), .A2(n_2372), .ZN(n_2400));
   XOR2_X1 i_1625 (.A(n_2400), .B(n_2374), .Z(n_2267));
   INV_X1 i_1626 (.A(n_2378), .ZN(n_2401));
   NAND2_X1 i_1627 (.A1(n_2401), .A2(n_2375), .ZN(n_2402));
   XOR2_X1 i_1628 (.A(n_2402), .B(n_2379), .Z(n_2274));
   INV_X1 i_1629 (.A(n_2381), .ZN(n_2403));
   NAND2_X1 i_1630 (.A1(n_2403), .A2(n_2380), .ZN(n_2405));
   XOR2_X1 i_1631 (.A(n_2405), .B(n_2382), .Z(n_2281));
   INV_X1 i_1632 (.A(n_2386), .ZN(n_2406));
   NAND2_X1 i_1633 (.A1(n_2406), .A2(n_2385), .ZN(n_2407));
   XOR2_X1 i_1634 (.A(n_2407), .B(n_2387), .Z(n_2288));
   INV_X1 i_1635 (.A(n_2389), .ZN(n_2408));
   NAND2_X1 i_1636 (.A1(n_2408), .A2(n_2388), .ZN(n_2409));
   XOR2_X1 i_1637 (.A(n_2409), .B(n_2392), .Z(n_2295));
   INV_X1 i_1638 (.A(n_712), .ZN(n_2410));
   NAND2_X1 i_1639 (.A1(n_2410), .A2(n_713), .ZN(n_2413));
   XOR2_X1 i_1640 (.A(n_2413), .B(n_711), .Z(n_2302));
   INV_X1 i_1641 (.A(n_709), .ZN(n_2414));
   NAND2_X1 i_1642 (.A1(n_2414), .A2(n_710), .ZN(n_2415));
   XOR2_X1 i_1643 (.A(n_2415), .B(n_708), .Z(n_2309));
   NAND4_X1 i_1644 (.A1(in1[23]), .A2(in1[22]), .A3(in2[2]), .A4(in2[1]), 
      .ZN(n_2416));
   AOI22_X1 i_1645 (.A1(in1[23]), .A2(in2[1]), .B1(in1[22]), .B2(in2[2]), 
      .ZN(n_2449));
   NAND2_X1 i_1646 (.A1(in1[21]), .A2(in2[3]), .ZN(n_2450));
   OAI21_X1 i_1647 (.A(n_2416), .B1(n_2449), .B2(n_2450), .ZN(n_2453));
   AOI21_X1 i_1648 (.A(n_2453), .B1(in1[25]), .B2(in2[0]), .ZN(n_2454));
   NAND2_X1 i_1649 (.A1(in1[24]), .A2(in2[1]), .ZN(n_2455));
   NAND3_X1 i_1650 (.A1(n_2453), .A2(in1[25]), .A3(in2[0]), .ZN(n_2456));
   AOI21_X1 i_1651 (.A(n_2454), .B1(n_2455), .B2(n_2456), .ZN(n_2215));
   NAND4_X1 i_1652 (.A1(in2[24]), .A2(in2[23]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2457));
   AOI22_X1 i_1653 (.A1(in2[23]), .A2(in1[2]), .B1(in2[24]), .B2(in1[1]), 
      .ZN(n_2460));
   NAND2_X1 i_1654 (.A1(in2[25]), .A2(in1[0]), .ZN(n_2461));
   OAI21_X1 i_1655 (.A(n_2457), .B1(n_2460), .B2(n_2461), .ZN(n_2160));
   NOR2_X1 i_1656 (.A1(n_3572), .A2(n_598), .ZN(n_2462));
   NAND3_X1 i_1657 (.A1(n_2462), .A2(in2[21]), .A3(in1[4]), .ZN(n_2463));
   AOI21_X1 i_1658 (.A(n_2462), .B1(in2[21]), .B2(in1[4]), .ZN(n_2464));
   NAND2_X1 i_1659 (.A1(in2[22]), .A2(in1[3]), .ZN(n_2467));
   OAI21_X1 i_1660 (.A(n_2463), .B1(n_2464), .B2(n_2467), .ZN(n_2167));
   NAND4_X1 i_1661 (.A1(in2[18]), .A2(in2[17]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2468));
   AOI22_X1 i_1662 (.A1(in2[17]), .A2(in1[8]), .B1(in2[18]), .B2(in1[7]), 
      .ZN(n_2469));
   NAND2_X1 i_1663 (.A1(in2[19]), .A2(in1[6]), .ZN(n_2470));
   OAI21_X1 i_1664 (.A(n_2468), .B1(n_2469), .B2(n_2470), .ZN(n_2174));
   NAND4_X1 i_1665 (.A1(in2[15]), .A2(in2[14]), .A3(in1[11]), .A4(in1[10]), 
      .ZN(n_2471));
   AOI22_X1 i_1666 (.A1(in2[14]), .A2(in1[11]), .B1(in2[15]), .B2(in1[10]), 
      .ZN(n_2474));
   NAND2_X1 i_1667 (.A1(in2[16]), .A2(in1[9]), .ZN(n_2475));
   OAI21_X1 i_1668 (.A(n_2471), .B1(n_2474), .B2(n_2475), .ZN(n_2181));
   NAND4_X1 i_1669 (.A1(in1[14]), .A2(in1[13]), .A3(in2[12]), .A4(in2[11]), 
      .ZN(n_2476));
   AOI22_X1 i_1670 (.A1(in1[14]), .A2(in2[11]), .B1(in1[13]), .B2(in2[12]), 
      .ZN(n_2477));
   NAND2_X1 i_1671 (.A1(in2[13]), .A2(in1[12]), .ZN(n_2478));
   OAI21_X1 i_1672 (.A(n_2476), .B1(n_2477), .B2(n_2478), .ZN(n_2188));
   NAND4_X1 i_1673 (.A1(in1[17]), .A2(in1[16]), .A3(in2[9]), .A4(in2[8]), 
      .ZN(n_2481));
   AOI22_X1 i_1674 (.A1(in1[17]), .A2(in2[8]), .B1(in1[16]), .B2(in2[9]), 
      .ZN(n_2482));
   NAND2_X1 i_1675 (.A1(in1[15]), .A2(in2[10]), .ZN(n_2483));
   OAI21_X1 i_1676 (.A(n_2481), .B1(n_2482), .B2(n_2483), .ZN(n_2195));
   NAND4_X1 i_1677 (.A1(in1[20]), .A2(in1[19]), .A3(in2[6]), .A4(in2[5]), 
      .ZN(n_2484));
   AOI22_X1 i_1678 (.A1(in1[20]), .A2(in2[5]), .B1(in1[19]), .B2(in2[6]), 
      .ZN(n_2485));
   NAND2_X1 i_1679 (.A1(in1[18]), .A2(in2[7]), .ZN(n_2488));
   OAI21_X1 i_1680 (.A(n_2484), .B1(n_2485), .B2(n_2488), .ZN(n_2202));
   NAND4_X1 i_1681 (.A1(in1[23]), .A2(in1[22]), .A3(in2[2]), .A4(in2[3]), 
      .ZN(n_2489));
   AOI22_X1 i_1682 (.A1(in1[23]), .A2(in2[2]), .B1(in1[22]), .B2(in2[3]), 
      .ZN(n_2490));
   NAND2_X1 i_1683 (.A1(in1[21]), .A2(in2[4]), .ZN(n_2491));
   OAI21_X1 i_1684 (.A(n_2489), .B1(n_2490), .B2(n_2491), .ZN(n_2209));
   INV_X1 i_1685 (.A(n_2460), .ZN(n_2492));
   NAND2_X1 i_1686 (.A1(n_2492), .A2(n_2457), .ZN(n_2495));
   XOR2_X1 i_1687 (.A(n_2495), .B(n_2461), .Z(n_2159));
   INV_X1 i_1688 (.A(n_2464), .ZN(n_2496));
   NAND2_X1 i_1689 (.A1(n_2463), .A2(n_2496), .ZN(n_2497));
   XOR2_X1 i_1690 (.A(n_2497), .B(n_2467), .Z(n_2166));
   INV_X1 i_1691 (.A(n_2469), .ZN(n_2498));
   NAND2_X1 i_1692 (.A1(n_2498), .A2(n_2468), .ZN(n_2499));
   XOR2_X1 i_1693 (.A(n_2499), .B(n_2470), .Z(n_2173));
   INV_X1 i_1694 (.A(n_2474), .ZN(n_2502));
   NAND2_X1 i_1695 (.A1(n_2502), .A2(n_2471), .ZN(n_2503));
   XOR2_X1 i_1696 (.A(n_2503), .B(n_2475), .Z(n_2180));
   INV_X1 i_1697 (.A(n_2477), .ZN(n_2504));
   NAND2_X1 i_1698 (.A1(n_2504), .A2(n_2476), .ZN(n_2505));
   XOR2_X1 i_1699 (.A(n_2505), .B(n_2478), .Z(n_2187));
   INV_X1 i_1700 (.A(n_2482), .ZN(n_2506));
   NAND2_X1 i_1701 (.A1(n_2506), .A2(n_2481), .ZN(n_2509));
   XOR2_X1 i_1702 (.A(n_2509), .B(n_2483), .Z(n_2194));
   INV_X1 i_1703 (.A(n_2485), .ZN(n_2510));
   NAND2_X1 i_1704 (.A1(n_2510), .A2(n_2484), .ZN(n_2511));
   XOR2_X1 i_1705 (.A(n_2511), .B(n_2488), .Z(n_2201));
   INV_X1 i_1706 (.A(n_2490), .ZN(n_2512));
   NAND2_X1 i_1707 (.A1(n_2512), .A2(n_2489), .ZN(n_2515));
   XOR2_X1 i_1708 (.A(n_2515), .B(n_2491), .Z(n_2208));
   INV_X1 i_1709 (.A(n_2454), .ZN(n_2516));
   NAND2_X1 i_1710 (.A1(n_2516), .A2(n_2456), .ZN(n_2517));
   XOR2_X1 i_1711 (.A(n_2517), .B(n_2455), .Z(n_2214));
   NAND4_X1 i_1712 (.A1(in1[20]), .A2(in1[19]), .A3(in2[3]), .A4(in2[4]), 
      .ZN(n_2518));
   AOI22_X1 i_1713 (.A1(in1[20]), .A2(in2[3]), .B1(in1[19]), .B2(in2[4]), 
      .ZN(n_2519));
   NAND2_X1 i_1714 (.A1(in1[18]), .A2(in2[5]), .ZN(n_2554));
   OAI21_X1 i_1715 (.A(n_2518), .B1(n_2519), .B2(n_2554), .ZN(n_2555));
   NAND4_X1 i_1716 (.A1(in1[23]), .A2(in1[22]), .A3(in2[1]), .A4(in2[0]), 
      .ZN(n_2558));
   AOI22_X1 i_1717 (.A1(in1[23]), .A2(in2[0]), .B1(in1[22]), .B2(in2[1]), 
      .ZN(n_2559));
   NAND2_X1 i_1718 (.A1(in1[21]), .A2(in2[2]), .ZN(n_2560));
   OAI21_X1 i_1719 (.A(n_2558), .B1(n_2559), .B2(n_2560), .ZN(n_2561));
   NOR2_X1 i_1720 (.A1(n_2555), .A2(n_2561), .ZN(n_2562));
   NAND2_X1 i_1721 (.A1(in1[24]), .A2(in2[0]), .ZN(n_2565));
   NAND2_X1 i_1722 (.A1(n_2555), .A2(n_2561), .ZN(n_2566));
   AOI21_X1 i_1723 (.A(n_2562), .B1(n_2565), .B2(n_2566), .ZN(n_2124));
   NAND4_X1 i_1724 (.A1(in2[23]), .A2(in2[22]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2567));
   AOI22_X1 i_1725 (.A1(in2[22]), .A2(in1[2]), .B1(in2[23]), .B2(in1[1]), 
      .ZN(n_2568));
   NAND2_X1 i_1726 (.A1(in2[24]), .A2(in1[0]), .ZN(n_2569));
   OAI21_X1 i_1727 (.A(n_2567), .B1(n_2568), .B2(n_2569), .ZN(n_2068));
   NAND3_X1 i_1728 (.A1(n_2462), .A2(in2[19]), .A3(in1[4]), .ZN(n_2572));
   AOI22_X1 i_1729 (.A1(in2[19]), .A2(in1[5]), .B1(in2[20]), .B2(in1[4]), 
      .ZN(n_2573));
   NAND2_X1 i_1730 (.A1(in2[21]), .A2(in1[3]), .ZN(n_2574));
   OAI21_X1 i_1731 (.A(n_2572), .B1(n_2573), .B2(n_2574), .ZN(n_2075));
   NAND4_X1 i_1732 (.A1(in2[17]), .A2(in2[16]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2575));
   AOI22_X1 i_1733 (.A1(in2[16]), .A2(in1[8]), .B1(in2[17]), .B2(in1[7]), 
      .ZN(n_2576));
   NAND2_X1 i_1734 (.A1(in2[18]), .A2(in1[6]), .ZN(n_2579));
   OAI21_X1 i_1735 (.A(n_2575), .B1(n_2576), .B2(n_2579), .ZN(n_2082));
   NAND4_X1 i_1736 (.A1(in2[14]), .A2(in2[13]), .A3(in1[11]), .A4(in1[10]), 
      .ZN(n_2580));
   AOI22_X1 i_1737 (.A1(in2[13]), .A2(in1[11]), .B1(in2[14]), .B2(in1[10]), 
      .ZN(n_2581));
   NAND2_X1 i_1738 (.A1(in2[15]), .A2(in1[9]), .ZN(n_2582));
   OAI21_X1 i_1739 (.A(n_2580), .B1(n_2581), .B2(n_2582), .ZN(n_2089));
   NAND4_X1 i_1740 (.A1(in1[14]), .A2(in1[13]), .A3(in2[11]), .A4(in2[10]), 
      .ZN(n_2583));
   AOI22_X1 i_1741 (.A1(in1[14]), .A2(in2[10]), .B1(in1[13]), .B2(in2[11]), 
      .ZN(n_2586));
   NAND2_X1 i_1742 (.A1(in1[12]), .A2(in2[12]), .ZN(n_2587));
   OAI21_X1 i_1743 (.A(n_2583), .B1(n_2586), .B2(n_2587), .ZN(n_2096));
   NAND4_X1 i_1744 (.A1(in1[17]), .A2(in1[16]), .A3(in2[8]), .A4(in2[7]), 
      .ZN(n_2588));
   AOI22_X1 i_1745 (.A1(in1[17]), .A2(in2[7]), .B1(in1[16]), .B2(in2[8]), 
      .ZN(n_2589));
   NAND2_X1 i_1746 (.A1(in1[15]), .A2(in2[9]), .ZN(n_2590));
   OAI21_X1 i_1747 (.A(n_2588), .B1(n_2589), .B2(n_2590), .ZN(n_2103));
   NAND4_X1 i_1748 (.A1(in1[20]), .A2(in1[19]), .A3(in2[4]), .A4(in2[5]), 
      .ZN(n_2593));
   AOI22_X1 i_1749 (.A1(in1[20]), .A2(in2[4]), .B1(in1[19]), .B2(in2[5]), 
      .ZN(n_2594));
   NAND2_X1 i_1750 (.A1(in1[18]), .A2(in2[6]), .ZN(n_2595));
   OAI21_X1 i_1751 (.A(n_2593), .B1(n_2594), .B2(n_2595), .ZN(n_2110));
   INV_X1 i_1752 (.A(n_2562), .ZN(n_2596));
   NAND2_X1 i_1753 (.A1(n_2596), .A2(n_2566), .ZN(n_2597));
   XOR2_X1 i_1754 (.A(n_2597), .B(n_2565), .Z(n_2123));
   INV_X1 i_1755 (.A(n_2568), .ZN(n_2600));
   NAND2_X1 i_1756 (.A1(n_2600), .A2(n_2567), .ZN(n_2601));
   XOR2_X1 i_1757 (.A(n_2601), .B(n_2569), .Z(n_2067));
   INV_X1 i_1758 (.A(n_2573), .ZN(n_2602));
   NAND2_X1 i_1759 (.A1(n_2572), .A2(n_2602), .ZN(n_2603));
   XOR2_X1 i_1760 (.A(n_2603), .B(n_2574), .Z(n_2074));
   INV_X1 i_1761 (.A(n_2576), .ZN(n_2604));
   NAND2_X1 i_1762 (.A1(n_2604), .A2(n_2575), .ZN(n_2607));
   XOR2_X1 i_1763 (.A(n_2607), .B(n_2579), .Z(n_2081));
   INV_X1 i_1764 (.A(n_2581), .ZN(n_2608));
   NAND2_X1 i_1765 (.A1(n_2608), .A2(n_2580), .ZN(n_2609));
   XOR2_X1 i_1766 (.A(n_2609), .B(n_2582), .Z(n_2088));
   INV_X1 i_1767 (.A(n_2586), .ZN(n_2610));
   NAND2_X1 i_1768 (.A1(n_2610), .A2(n_2583), .ZN(n_2611));
   XOR2_X1 i_1769 (.A(n_2611), .B(n_2587), .Z(n_2095));
   INV_X1 i_1770 (.A(n_2589), .ZN(n_2613));
   NAND2_X1 i_1771 (.A1(n_2613), .A2(n_2588), .ZN(n_2614));
   XOR2_X1 i_1772 (.A(n_2614), .B(n_2590), .Z(n_2102));
   INV_X1 i_1773 (.A(n_2594), .ZN(n_2615));
   NAND2_X1 i_1774 (.A1(n_2615), .A2(n_2593), .ZN(n_2616));
   XOR2_X1 i_1775 (.A(n_2616), .B(n_2595), .Z(n_2109));
   INV_X1 i_1776 (.A(n_2449), .ZN(n_2617));
   NAND2_X1 i_1777 (.A1(n_2617), .A2(n_2416), .ZN(n_2618));
   XOR2_X1 i_1778 (.A(n_2618), .B(n_2450), .Z(n_2116));
   NAND4_X1 i_1779 (.A1(in2[22]), .A2(in2[21]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2620));
   AOI22_X1 i_1780 (.A1(in2[21]), .A2(in1[2]), .B1(in2[22]), .B2(in1[1]), 
      .ZN(n_2621));
   NAND2_X1 i_1781 (.A1(in2[23]), .A2(in1[0]), .ZN(n_2622));
   OAI21_X1 i_1782 (.A(n_2620), .B1(n_2621), .B2(n_2622), .ZN(n_1984));
   NOR2_X1 i_1783 (.A1(n_2859), .A2(n_598), .ZN(n_2623));
   NAND3_X1 i_1784 (.A1(n_2623), .A2(in2[19]), .A3(in1[4]), .ZN(n_2660));
   AOI21_X1 i_1785 (.A(n_2623), .B1(in2[19]), .B2(in1[4]), .ZN(n_2661));
   NAND2_X1 i_1786 (.A1(in2[20]), .A2(in1[3]), .ZN(n_2664));
   OAI21_X1 i_1787 (.A(n_2660), .B1(n_2661), .B2(n_2664), .ZN(n_1991));
   NAND4_X1 i_1788 (.A1(in2[16]), .A2(in2[15]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2665));
   AOI22_X1 i_1789 (.A1(in2[15]), .A2(in1[8]), .B1(in2[16]), .B2(in1[7]), 
      .ZN(n_2666));
   NAND2_X1 i_1790 (.A1(in2[17]), .A2(in1[6]), .ZN(n_2667));
   OAI21_X1 i_1791 (.A(n_2665), .B1(n_2666), .B2(n_2667), .ZN(n_1998));
   NAND4_X1 i_1792 (.A1(in2[13]), .A2(in1[11]), .A3(in2[12]), .A4(in1[10]), 
      .ZN(n_2668));
   AOI22_X1 i_1793 (.A1(in1[11]), .A2(in2[12]), .B1(in2[13]), .B2(in1[10]), 
      .ZN(n_2671));
   NAND2_X1 i_1794 (.A1(in2[14]), .A2(in1[9]), .ZN(n_2672));
   OAI21_X1 i_1795 (.A(n_2668), .B1(n_2671), .B2(n_2672), .ZN(n_2005));
   NAND4_X1 i_1796 (.A1(in1[14]), .A2(in1[13]), .A3(in2[10]), .A4(in2[9]), 
      .ZN(n_2673));
   AOI22_X1 i_1797 (.A1(in1[14]), .A2(in2[9]), .B1(in1[13]), .B2(in2[10]), 
      .ZN(n_2674));
   NAND2_X1 i_1798 (.A1(in1[12]), .A2(in2[11]), .ZN(n_2675));
   OAI21_X1 i_1799 (.A(n_2673), .B1(n_2674), .B2(n_2675), .ZN(n_2012));
   NAND4_X1 i_1800 (.A1(in1[17]), .A2(in1[16]), .A3(in2[7]), .A4(in2[6]), 
      .ZN(n_2678));
   AOI22_X1 i_1801 (.A1(in1[17]), .A2(in2[6]), .B1(in1[16]), .B2(in2[7]), 
      .ZN(n_2679));
   NAND2_X1 i_1802 (.A1(in1[15]), .A2(in2[8]), .ZN(n_2680));
   OAI21_X1 i_1803 (.A(n_2678), .B1(n_2679), .B2(n_2680), .ZN(n_2019));
   INV_X1 i_1804 (.A(n_2621), .ZN(n_2681));
   NAND2_X1 i_1805 (.A1(n_2681), .A2(n_2620), .ZN(n_2682));
   XOR2_X1 i_1806 (.A(n_2682), .B(n_2622), .Z(n_1983));
   INV_X1 i_1807 (.A(n_2661), .ZN(n_2685));
   NAND2_X1 i_1808 (.A1(n_2660), .A2(n_2685), .ZN(n_2686));
   XOR2_X1 i_1809 (.A(n_2686), .B(n_2664), .Z(n_1990));
   INV_X1 i_1810 (.A(n_2666), .ZN(n_2687));
   NAND2_X1 i_1811 (.A1(n_2687), .A2(n_2665), .ZN(n_2688));
   XOR2_X1 i_1812 (.A(n_2688), .B(n_2667), .Z(n_1997));
   INV_X1 i_1813 (.A(n_2671), .ZN(n_2689));
   NAND2_X1 i_1814 (.A1(n_2689), .A2(n_2668), .ZN(n_2692));
   XOR2_X1 i_1815 (.A(n_2692), .B(n_2672), .Z(n_2004));
   INV_X1 i_1816 (.A(n_2674), .ZN(n_2693));
   NAND2_X1 i_1817 (.A1(n_2693), .A2(n_2673), .ZN(n_2694));
   XOR2_X1 i_1818 (.A(n_2694), .B(n_2675), .Z(n_2011));
   INV_X1 i_1819 (.A(n_2679), .ZN(n_2695));
   NAND2_X1 i_1820 (.A1(n_2695), .A2(n_2678), .ZN(n_2696));
   XOR2_X1 i_1821 (.A(n_2696), .B(n_2680), .Z(n_2018));
   INV_X1 i_1822 (.A(n_2519), .ZN(n_2699));
   NAND2_X1 i_1823 (.A1(n_2699), .A2(n_2518), .ZN(n_2700));
   XOR2_X1 i_1824 (.A(n_2700), .B(n_2554), .Z(n_2025));
   INV_X1 i_1825 (.A(n_2559), .ZN(n_2701));
   NAND2_X1 i_1826 (.A1(n_2701), .A2(n_2558), .ZN(n_2702));
   XOR2_X1 i_1827 (.A(n_2702), .B(n_2560), .Z(n_2032));
   NAND4_X1 i_1828 (.A1(in1[20]), .A2(in1[19]), .A3(in2[2]), .A4(in2[1]), 
      .ZN(n_2703));
   AOI22_X1 i_1829 (.A1(in1[20]), .A2(in2[1]), .B1(in1[19]), .B2(in2[2]), 
      .ZN(n_2706));
   NAND2_X1 i_1830 (.A1(in1[18]), .A2(in2[3]), .ZN(n_2707));
   OAI21_X1 i_1831 (.A(n_2703), .B1(n_2706), .B2(n_2707), .ZN(n_2708));
   AOI21_X1 i_1832 (.A(n_2708), .B1(in1[22]), .B2(in2[0]), .ZN(n_2709));
   NAND2_X1 i_1833 (.A1(in1[21]), .A2(in2[1]), .ZN(n_2710));
   NAND3_X1 i_1834 (.A1(n_2708), .A2(in1[22]), .A3(in2[0]), .ZN(n_2713));
   AOI21_X1 i_1835 (.A(n_2709), .B1(n_2710), .B2(n_2713), .ZN(n_1949));
   NAND4_X1 i_1836 (.A1(in2[21]), .A2(in2[20]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2714));
   AOI22_X1 i_1837 (.A1(in2[20]), .A2(in1[2]), .B1(in2[21]), .B2(in1[1]), 
      .ZN(n_2715));
   NAND2_X1 i_1838 (.A1(in2[22]), .A2(in1[0]), .ZN(n_2716));
   OAI21_X1 i_1839 (.A(n_2714), .B1(n_2715), .B2(n_2716), .ZN(n_1901));
   NOR2_X1 i_1840 (.A1(n_2857), .A2(n_598), .ZN(n_2717));
   NAND3_X1 i_1841 (.A1(n_2717), .A2(in2[18]), .A3(in1[4]), .ZN(n_2720));
   AOI21_X1 i_1842 (.A(n_2717), .B1(in2[18]), .B2(in1[4]), .ZN(n_2721));
   NAND2_X1 i_1843 (.A1(in2[19]), .A2(in1[3]), .ZN(n_2722));
   OAI21_X1 i_1844 (.A(n_2720), .B1(n_2721), .B2(n_2722), .ZN(n_1908));
   NAND4_X1 i_1845 (.A1(in2[15]), .A2(in2[14]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2723));
   AOI22_X1 i_1846 (.A1(in2[14]), .A2(in1[8]), .B1(in2[15]), .B2(in1[7]), 
      .ZN(n_2724));
   NAND2_X1 i_1847 (.A1(in2[16]), .A2(in1[6]), .ZN(n_2726));
   OAI21_X1 i_1848 (.A(n_2723), .B1(n_2724), .B2(n_2726), .ZN(n_1915));
   NAND4_X1 i_1849 (.A1(in1[11]), .A2(in2[12]), .A3(in2[11]), .A4(in1[10]), 
      .ZN(n_2727));
   AOI22_X1 i_1850 (.A1(in1[11]), .A2(in2[11]), .B1(in2[12]), .B2(in1[10]), 
      .ZN(n_2728));
   NAND2_X1 i_1851 (.A1(in2[13]), .A2(in1[9]), .ZN(n_2729));
   OAI21_X1 i_1852 (.A(n_2727), .B1(n_2728), .B2(n_2729), .ZN(n_1922));
   NAND4_X1 i_1853 (.A1(in1[14]), .A2(in1[13]), .A3(in2[9]), .A4(in2[8]), 
      .ZN(n_2730));
   AOI22_X1 i_1854 (.A1(in1[14]), .A2(in2[8]), .B1(in1[13]), .B2(in2[9]), 
      .ZN(n_2731));
   NAND2_X1 i_1855 (.A1(in1[12]), .A2(in2[10]), .ZN(n_2734));
   OAI21_X1 i_1856 (.A(n_2730), .B1(n_2731), .B2(n_2734), .ZN(n_1929));
   NAND4_X1 i_1857 (.A1(in1[17]), .A2(in1[16]), .A3(in2[6]), .A4(in2[5]), 
      .ZN(n_2735));
   AOI22_X1 i_1858 (.A1(in1[17]), .A2(in2[5]), .B1(in1[16]), .B2(in2[6]), 
      .ZN(n_2736));
   NAND2_X1 i_1859 (.A1(in1[15]), .A2(in2[7]), .ZN(n_2737));
   OAI21_X1 i_1860 (.A(n_2735), .B1(n_2736), .B2(n_2737), .ZN(n_1936));
   NAND4_X1 i_1861 (.A1(in1[20]), .A2(in1[19]), .A3(in2[2]), .A4(in2[3]), 
      .ZN(n_2774));
   AOI22_X1 i_1862 (.A1(in1[20]), .A2(in2[2]), .B1(in1[19]), .B2(in2[3]), 
      .ZN(n_2777));
   NAND2_X1 i_1863 (.A1(in1[18]), .A2(in2[4]), .ZN(n_2778));
   OAI21_X1 i_1864 (.A(n_2774), .B1(n_2777), .B2(n_2778), .ZN(n_1943));
   INV_X1 i_1865 (.A(n_2715), .ZN(n_2779));
   NAND2_X1 i_1866 (.A1(n_2779), .A2(n_2714), .ZN(n_2780));
   XOR2_X1 i_1867 (.A(n_2780), .B(n_2716), .Z(n_1900));
   INV_X1 i_1868 (.A(n_2721), .ZN(n_2781));
   NAND2_X1 i_1869 (.A1(n_2720), .A2(n_2781), .ZN(n_2782));
   XOR2_X1 i_1870 (.A(n_2782), .B(n_2722), .Z(n_1907));
   INV_X1 i_1871 (.A(n_2724), .ZN(n_2783));
   NAND2_X1 i_1872 (.A1(n_2783), .A2(n_2723), .ZN(n_2786));
   XOR2_X1 i_1873 (.A(n_2786), .B(n_2726), .Z(n_1914));
   INV_X1 i_1874 (.A(n_2728), .ZN(n_2787));
   NAND2_X1 i_1875 (.A1(n_2787), .A2(n_2727), .ZN(n_2788));
   XOR2_X1 i_1876 (.A(n_2788), .B(n_2729), .Z(n_1921));
   INV_X1 i_1877 (.A(n_2731), .ZN(n_2789));
   NAND2_X1 i_1878 (.A1(n_2789), .A2(n_2730), .ZN(n_2790));
   XOR2_X1 i_1879 (.A(n_2790), .B(n_2734), .Z(n_1928));
   INV_X1 i_1880 (.A(n_2736), .ZN(n_2793));
   NAND2_X1 i_1881 (.A1(n_2793), .A2(n_2735), .ZN(n_2794));
   XOR2_X1 i_1882 (.A(n_2794), .B(n_2737), .Z(n_1935));
   INV_X1 i_1883 (.A(n_2777), .ZN(n_2795));
   NAND2_X1 i_1884 (.A1(n_2795), .A2(n_2774), .ZN(n_2796));
   XOR2_X1 i_1885 (.A(n_2796), .B(n_2778), .Z(n_1942));
   INV_X1 i_1886 (.A(n_2709), .ZN(n_2797));
   NAND2_X1 i_1887 (.A1(n_2797), .A2(n_2713), .ZN(n_2800));
   XOR2_X1 i_1888 (.A(n_2800), .B(n_2710), .Z(n_1948));
   NAND4_X1 i_1889 (.A1(in1[17]), .A2(in1[16]), .A3(in2[3]), .A4(in2[4]), 
      .ZN(n_2801));
   AOI22_X1 i_1890 (.A1(in1[17]), .A2(in2[3]), .B1(in1[16]), .B2(in2[4]), 
      .ZN(n_2802));
   NAND2_X1 i_1891 (.A1(in1[15]), .A2(in2[5]), .ZN(n_2803));
   OAI21_X1 i_1892 (.A(n_2801), .B1(n_2802), .B2(n_2803), .ZN(n_2804));
   NAND4_X1 i_1893 (.A1(in1[20]), .A2(in1[19]), .A3(in2[1]), .A4(in2[0]), 
      .ZN(n_2807));
   AOI22_X1 i_1894 (.A1(in1[20]), .A2(in2[0]), .B1(in1[19]), .B2(in2[1]), 
      .ZN(n_2808));
   NAND2_X1 i_1895 (.A1(in1[18]), .A2(in2[2]), .ZN(n_2809));
   OAI21_X1 i_1896 (.A(n_2807), .B1(n_2808), .B2(n_2809), .ZN(n_2810));
   NOR2_X1 i_1897 (.A1(n_2804), .A2(n_2810), .ZN(n_2811));
   NAND2_X1 i_1898 (.A1(in1[21]), .A2(in2[0]), .ZN(n_2814));
   NAND2_X1 i_1899 (.A1(n_2804), .A2(n_2810), .ZN(n_2815));
   AOI21_X1 i_1900 (.A(n_2811), .B1(n_2814), .B2(n_2815), .ZN(n_1869));
   NAND4_X1 i_1901 (.A1(in2[20]), .A2(in2[19]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2816));
   AOI22_X1 i_1902 (.A1(in2[19]), .A2(in1[2]), .B1(in2[20]), .B2(in1[1]), 
      .ZN(n_2817));
   NAND2_X1 i_1903 (.A1(in2[21]), .A2(in1[0]), .ZN(n_2818));
   OAI21_X1 i_1904 (.A(n_2816), .B1(n_2817), .B2(n_2818), .ZN(n_1820));
   NAND3_X1 i_1905 (.A1(n_2717), .A2(in2[16]), .A3(in1[4]), .ZN(n_2821));
   AOI22_X1 i_1906 (.A1(in2[16]), .A2(in1[5]), .B1(in2[17]), .B2(in1[4]), 
      .ZN(n_2822));
   NAND2_X1 i_1907 (.A1(in2[18]), .A2(in1[3]), .ZN(n_2823));
   OAI21_X1 i_1908 (.A(n_2821), .B1(n_2822), .B2(n_2823), .ZN(n_1827));
   NAND4_X1 i_1909 (.A1(in2[14]), .A2(in2[13]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2824));
   AOI22_X1 i_1910 (.A1(in2[13]), .A2(in1[8]), .B1(in2[14]), .B2(in1[7]), 
      .ZN(n_2825));
   NAND2_X1 i_1911 (.A1(in2[15]), .A2(in1[6]), .ZN(n_2828));
   OAI21_X1 i_1912 (.A(n_2824), .B1(n_2825), .B2(n_2828), .ZN(n_1834));
   NAND4_X1 i_1913 (.A1(in1[11]), .A2(in2[11]), .A3(in1[10]), .A4(in2[10]), 
      .ZN(n_2829));
   AOI22_X1 i_1914 (.A1(in1[11]), .A2(in2[10]), .B1(in2[11]), .B2(in1[10]), 
      .ZN(n_2830));
   NAND2_X1 i_1915 (.A1(in2[12]), .A2(in1[9]), .ZN(n_2831));
   OAI21_X1 i_1916 (.A(n_2829), .B1(n_2830), .B2(n_2831), .ZN(n_1841));
   NAND4_X1 i_1917 (.A1(in1[14]), .A2(in1[13]), .A3(in2[8]), .A4(in2[7]), 
      .ZN(n_2832));
   AOI22_X1 i_1918 (.A1(in1[14]), .A2(in2[7]), .B1(in1[13]), .B2(in2[8]), 
      .ZN(n_2835));
   NAND2_X1 i_1919 (.A1(in1[12]), .A2(in2[9]), .ZN(n_2836));
   OAI21_X1 i_1920 (.A(n_2832), .B1(n_2835), .B2(n_2836), .ZN(n_1848));
   NAND4_X1 i_1921 (.A1(in1[17]), .A2(in1[16]), .A3(in2[4]), .A4(in2[5]), 
      .ZN(n_2837));
   AOI22_X1 i_1922 (.A1(in1[17]), .A2(in2[4]), .B1(in1[16]), .B2(in2[5]), 
      .ZN(n_2838));
   NAND2_X1 i_1923 (.A1(in1[15]), .A2(in2[6]), .ZN(n_2839));
   OAI21_X1 i_1924 (.A(n_2837), .B1(n_2838), .B2(n_2839), .ZN(n_1855));
   INV_X1 i_1925 (.A(n_2811), .ZN(n_2841));
   NAND2_X1 i_1926 (.A1(n_2841), .A2(n_2815), .ZN(n_2842));
   XOR2_X1 i_1927 (.A(n_2842), .B(n_2814), .Z(n_1868));
   INV_X1 i_1928 (.A(n_2817), .ZN(n_2843));
   NAND2_X1 i_1929 (.A1(n_2843), .A2(n_2816), .ZN(n_2844));
   XOR2_X1 i_1930 (.A(n_2844), .B(n_2818), .Z(n_1819));
   INV_X1 i_1931 (.A(n_2822), .ZN(n_2845));
   NAND2_X1 i_1932 (.A1(n_2821), .A2(n_2845), .ZN(n_2846));
   XOR2_X1 i_1933 (.A(n_2846), .B(n_2823), .Z(n_1826));
   INV_X1 i_1934 (.A(n_2825), .ZN(n_2849));
   NAND2_X1 i_1935 (.A1(n_2849), .A2(n_2824), .ZN(n_2850));
   XOR2_X1 i_1936 (.A(n_2850), .B(n_2828), .Z(n_1833));
   INV_X1 i_1937 (.A(n_2830), .ZN(n_2851));
   NAND2_X1 i_1938 (.A1(n_2851), .A2(n_2829), .ZN(n_2852));
   XOR2_X1 i_1939 (.A(n_2852), .B(n_2831), .Z(n_1840));
   INV_X1 i_1940 (.A(n_2835), .ZN(n_2891));
   NAND2_X1 i_1941 (.A1(n_2891), .A2(n_2832), .ZN(n_2894));
   XOR2_X1 i_1942 (.A(n_2894), .B(n_2836), .Z(n_1847));
   INV_X1 i_1943 (.A(n_2838), .ZN(n_2895));
   NAND2_X1 i_1944 (.A1(n_2895), .A2(n_2837), .ZN(n_2896));
   XOR2_X1 i_1945 (.A(n_2896), .B(n_2839), .Z(n_1854));
   INV_X1 i_1946 (.A(n_2706), .ZN(n_2899));
   NAND2_X1 i_1947 (.A1(n_2899), .A2(n_2703), .ZN(n_2900));
   XOR2_X1 i_1948 (.A(n_2900), .B(n_2707), .Z(n_1861));
   NAND4_X1 i_1949 (.A1(in2[19]), .A2(in2[18]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2901));
   AOI22_X1 i_1950 (.A1(in2[18]), .A2(in1[2]), .B1(in2[19]), .B2(in1[1]), 
      .ZN(n_2902));
   NAND2_X1 i_1951 (.A1(in2[20]), .A2(in1[0]), .ZN(n_2903));
   OAI21_X1 i_1952 (.A(n_2901), .B1(n_2902), .B2(n_2903), .ZN(n_1747));
   NOR2_X1 i_1953 (.A1(n_790), .A2(n_598), .ZN(n_2906));
   NAND3_X1 i_1954 (.A1(n_2906), .A2(in2[16]), .A3(in1[4]), .ZN(n_2907));
   AOI21_X1 i_1955 (.A(n_2906), .B1(in2[16]), .B2(in1[4]), .ZN(n_2908));
   NAND2_X1 i_1956 (.A1(in2[17]), .A2(in1[3]), .ZN(n_2909));
   OAI21_X1 i_1957 (.A(n_2907), .B1(n_2908), .B2(n_2909), .ZN(n_1754));
   NAND4_X1 i_1958 (.A1(in2[13]), .A2(in2[12]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2910));
   AOI22_X1 i_1959 (.A1(in2[12]), .A2(in1[8]), .B1(in2[13]), .B2(in1[7]), 
      .ZN(n_2913));
   NAND2_X1 i_1960 (.A1(in2[14]), .A2(in1[6]), .ZN(n_2914));
   OAI21_X1 i_1961 (.A(n_2910), .B1(n_2913), .B2(n_2914), .ZN(n_1761));
   NAND4_X1 i_1962 (.A1(in1[11]), .A2(in1[10]), .A3(in2[10]), .A4(in2[9]), 
      .ZN(n_2915));
   AOI22_X1 i_1963 (.A1(in1[11]), .A2(in2[9]), .B1(in1[10]), .B2(in2[10]), 
      .ZN(n_2916));
   NAND2_X1 i_1964 (.A1(in2[11]), .A2(in1[9]), .ZN(n_2917));
   OAI21_X1 i_1965 (.A(n_2915), .B1(n_2916), .B2(n_2917), .ZN(n_1768));
   NAND4_X1 i_1966 (.A1(in1[14]), .A2(in1[13]), .A3(in2[7]), .A4(in2[6]), 
      .ZN(n_2920));
   AOI22_X1 i_1967 (.A1(in1[14]), .A2(in2[6]), .B1(in1[13]), .B2(in2[7]), 
      .ZN(n_2921));
   NAND2_X1 i_1968 (.A1(in1[12]), .A2(in2[8]), .ZN(n_2922));
   OAI21_X1 i_1969 (.A(n_2920), .B1(n_2921), .B2(n_2922), .ZN(n_1775));
   INV_X1 i_1970 (.A(n_2902), .ZN(n_2923));
   NAND2_X1 i_1971 (.A1(n_2923), .A2(n_2901), .ZN(n_2924));
   XOR2_X1 i_1972 (.A(n_2924), .B(n_2903), .Z(n_1746));
   INV_X1 i_1973 (.A(n_2908), .ZN(n_2927));
   NAND2_X1 i_1974 (.A1(n_2907), .A2(n_2927), .ZN(n_2928));
   XOR2_X1 i_1975 (.A(n_2928), .B(n_2909), .Z(n_1753));
   INV_X1 i_1976 (.A(n_2913), .ZN(n_2929));
   NAND2_X1 i_1977 (.A1(n_2929), .A2(n_2910), .ZN(n_2930));
   XOR2_X1 i_1978 (.A(n_2930), .B(n_2914), .Z(n_1760));
   INV_X1 i_1979 (.A(n_2916), .ZN(n_2931));
   NAND2_X1 i_1980 (.A1(n_2931), .A2(n_2915), .ZN(n_2934));
   XOR2_X1 i_1981 (.A(n_2934), .B(n_2917), .Z(n_1767));
   INV_X1 i_1982 (.A(n_2921), .ZN(n_2935));
   NAND2_X1 i_1983 (.A1(n_2935), .A2(n_2920), .ZN(n_2936));
   XOR2_X1 i_1984 (.A(n_2936), .B(n_2922), .Z(n_1774));
   INV_X1 i_1985 (.A(n_2802), .ZN(n_2937));
   NAND2_X1 i_1986 (.A1(n_2937), .A2(n_2801), .ZN(n_2938));
   XOR2_X1 i_1987 (.A(n_2938), .B(n_2803), .Z(n_1781));
   INV_X1 i_1988 (.A(n_2808), .ZN(n_2941));
   NAND2_X1 i_1989 (.A1(n_2941), .A2(n_2807), .ZN(n_2942));
   XOR2_X1 i_1990 (.A(n_2942), .B(n_2809), .Z(n_1788));
   NAND4_X1 i_1991 (.A1(in1[17]), .A2(in1[16]), .A3(in2[2]), .A4(in2[1]), 
      .ZN(n_2943));
   AOI22_X1 i_1992 (.A1(in1[17]), .A2(in2[1]), .B1(in1[16]), .B2(in2[2]), 
      .ZN(n_2944));
   NAND2_X1 i_1993 (.A1(in1[15]), .A2(in2[3]), .ZN(n_2945));
   OAI21_X1 i_1994 (.A(n_2943), .B1(n_2944), .B2(n_2945), .ZN(n_2948));
   AOI21_X1 i_1995 (.A(n_2948), .B1(in1[19]), .B2(in2[0]), .ZN(n_2949));
   NAND2_X1 i_1996 (.A1(in1[18]), .A2(in2[1]), .ZN(n_2950));
   NAND3_X1 i_1997 (.A1(n_2948), .A2(in1[19]), .A3(in2[0]), .ZN(n_2951));
   AOI21_X1 i_1998 (.A(n_2949), .B1(n_2950), .B2(n_2951), .ZN(n_1716));
   NAND4_X1 i_1999 (.A1(in2[18]), .A2(in2[17]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_2952));
   AOI22_X1 i_2000 (.A1(in2[17]), .A2(in1[2]), .B1(in2[18]), .B2(in1[1]), 
      .ZN(n_2955));
   NAND2_X1 i_2001 (.A1(in2[19]), .A2(in1[0]), .ZN(n_2956));
   OAI21_X1 i_2002 (.A(n_2952), .B1(n_2955), .B2(n_2956), .ZN(n_1675));
   NOR2_X1 i_2003 (.A1(n_788), .A2(n_598), .ZN(n_2957));
   NAND3_X1 i_2004 (.A1(n_2957), .A2(in2[15]), .A3(in1[4]), .ZN(n_2958));
   AOI21_X1 i_2005 (.A(n_2957), .B1(in2[15]), .B2(in1[4]), .ZN(n_2959));
   NAND2_X1 i_2006 (.A1(in2[16]), .A2(in1[3]), .ZN(n_2962));
   OAI21_X1 i_2007 (.A(n_2958), .B1(n_2959), .B2(n_2962), .ZN(n_1682));
   NAND4_X1 i_2008 (.A1(in2[12]), .A2(in2[11]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_2963));
   AOI22_X1 i_2009 (.A1(in2[11]), .A2(in1[8]), .B1(in2[12]), .B2(in1[7]), 
      .ZN(n_2964));
   NAND2_X1 i_2010 (.A1(in2[13]), .A2(in1[6]), .ZN(n_2965));
   OAI21_X1 i_2011 (.A(n_2963), .B1(n_2964), .B2(n_2965), .ZN(n_1689));
   NAND4_X1 i_2012 (.A1(in1[11]), .A2(in1[10]), .A3(in2[9]), .A4(in2[8]), 
      .ZN(n_3004));
   AOI22_X1 i_2013 (.A1(in1[11]), .A2(in2[8]), .B1(in1[10]), .B2(in2[9]), 
      .ZN(n_3007));
   NAND2_X1 i_2014 (.A1(in2[10]), .A2(in1[9]), .ZN(n_3008));
   OAI21_X1 i_2015 (.A(n_3004), .B1(n_3007), .B2(n_3008), .ZN(n_1696));
   NAND4_X1 i_2016 (.A1(in1[14]), .A2(in1[13]), .A3(in2[6]), .A4(in2[5]), 
      .ZN(n_3009));
   AOI22_X1 i_2017 (.A1(in1[14]), .A2(in2[5]), .B1(in1[13]), .B2(in2[6]), 
      .ZN(n_3010));
   NAND2_X1 i_2018 (.A1(in1[12]), .A2(in2[7]), .ZN(n_3011));
   OAI21_X1 i_2019 (.A(n_3009), .B1(n_3010), .B2(n_3011), .ZN(n_1703));
   NAND4_X1 i_2020 (.A1(in1[17]), .A2(in1[16]), .A3(in2[2]), .A4(in2[3]), 
      .ZN(n_3012));
   AOI22_X1 i_2021 (.A1(in1[17]), .A2(in2[2]), .B1(in1[16]), .B2(in2[3]), 
      .ZN(n_3013));
   NAND2_X1 i_2022 (.A1(in1[15]), .A2(in2[4]), .ZN(n_3016));
   OAI21_X1 i_2023 (.A(n_3012), .B1(n_3013), .B2(n_3016), .ZN(n_1710));
   INV_X1 i_2024 (.A(n_2955), .ZN(n_3017));
   NAND2_X1 i_2025 (.A1(n_3017), .A2(n_2952), .ZN(n_3018));
   XOR2_X1 i_2026 (.A(n_3018), .B(n_2956), .Z(n_1674));
   INV_X1 i_2027 (.A(n_2959), .ZN(n_3019));
   NAND2_X1 i_2028 (.A1(n_2958), .A2(n_3019), .ZN(n_3020));
   XOR2_X1 i_2029 (.A(n_3020), .B(n_2962), .Z(n_1681));
   INV_X1 i_2030 (.A(n_2964), .ZN(n_3023));
   NAND2_X1 i_2031 (.A1(n_3023), .A2(n_2963), .ZN(n_3024));
   XOR2_X1 i_2032 (.A(n_3024), .B(n_2965), .Z(n_1688));
   INV_X1 i_2033 (.A(n_3007), .ZN(n_3025));
   NAND2_X1 i_2034 (.A1(n_3025), .A2(n_3004), .ZN(n_3026));
   XOR2_X1 i_2035 (.A(n_3026), .B(n_3008), .Z(n_1695));
   INV_X1 i_2036 (.A(n_3010), .ZN(n_3027));
   NAND2_X1 i_2037 (.A1(n_3027), .A2(n_3009), .ZN(n_3030));
   XOR2_X1 i_2038 (.A(n_3030), .B(n_3011), .Z(n_1702));
   INV_X1 i_2039 (.A(n_3013), .ZN(n_3031));
   NAND2_X1 i_2040 (.A1(n_3031), .A2(n_3012), .ZN(n_3032));
   XOR2_X1 i_2041 (.A(n_3032), .B(n_3016), .Z(n_1709));
   INV_X1 i_2042 (.A(n_2949), .ZN(n_3033));
   NAND2_X1 i_2043 (.A1(n_3033), .A2(n_2951), .ZN(n_3034));
   XOR2_X1 i_2044 (.A(n_3034), .B(n_2950), .Z(n_1715));
   NAND4_X1 i_2045 (.A1(in1[14]), .A2(in1[13]), .A3(in2[3]), .A4(in2[4]), 
      .ZN(n_3037));
   AOI22_X1 i_2046 (.A1(in1[14]), .A2(in2[3]), .B1(in1[13]), .B2(in2[4]), 
      .ZN(n_3038));
   NAND2_X1 i_2047 (.A1(in1[12]), .A2(in2[5]), .ZN(n_3039));
   OAI21_X1 i_2048 (.A(n_3037), .B1(n_3038), .B2(n_3039), .ZN(n_3040));
   NAND4_X1 i_2049 (.A1(in1[17]), .A2(in1[16]), .A3(in2[1]), .A4(in2[0]), 
      .ZN(n_3041));
   AOI22_X1 i_2050 (.A1(in1[17]), .A2(in2[0]), .B1(in1[16]), .B2(in2[1]), 
      .ZN(n_3044));
   NAND2_X1 i_2051 (.A1(in1[15]), .A2(in2[2]), .ZN(n_3045));
   OAI21_X1 i_2052 (.A(n_3041), .B1(n_3044), .B2(n_3045), .ZN(n_3046));
   NOR2_X1 i_2053 (.A1(n_3040), .A2(n_3046), .ZN(n_3047));
   NAND2_X1 i_2054 (.A1(in1[18]), .A2(in2[0]), .ZN(n_3048));
   NAND2_X1 i_2055 (.A1(n_3040), .A2(n_3046), .ZN(n_3051));
   AOI21_X1 i_2056 (.A(n_3047), .B1(n_3048), .B2(n_3051), .ZN(n_1647));
   NAND4_X1 i_2057 (.A1(in2[17]), .A2(in2[16]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3052));
   AOI22_X1 i_2058 (.A1(in2[16]), .A2(in1[2]), .B1(in2[17]), .B2(in1[1]), 
      .ZN(n_3053));
   NAND2_X1 i_2059 (.A1(in2[18]), .A2(in1[0]), .ZN(n_3054));
   OAI21_X1 i_2060 (.A(n_3052), .B1(n_3053), .B2(n_3054), .ZN(n_1605));
   NAND3_X1 i_2061 (.A1(n_2957), .A2(in2[13]), .A3(in1[4]), .ZN(n_3055));
   AOI22_X1 i_2062 (.A1(in2[13]), .A2(in1[5]), .B1(in2[14]), .B2(in1[4]), 
      .ZN(n_3058));
   NAND2_X1 i_2063 (.A1(in2[15]), .A2(in1[3]), .ZN(n_3059));
   OAI21_X1 i_2064 (.A(n_3055), .B1(n_3058), .B2(n_3059), .ZN(n_1612));
   NAND4_X1 i_2065 (.A1(in2[11]), .A2(in2[10]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_3060));
   AOI22_X1 i_2066 (.A1(in2[10]), .A2(in1[8]), .B1(in2[11]), .B2(in1[7]), 
      .ZN(n_3061));
   NAND2_X1 i_2067 (.A1(in2[12]), .A2(in1[6]), .ZN(n_3062));
   OAI21_X1 i_2068 (.A(n_3060), .B1(n_3061), .B2(n_3062), .ZN(n_1619));
   NAND4_X1 i_2069 (.A1(in1[11]), .A2(in1[10]), .A3(in2[8]), .A4(in2[7]), 
      .ZN(n_3065));
   AOI22_X1 i_2070 (.A1(in1[11]), .A2(in2[7]), .B1(in1[10]), .B2(in2[8]), 
      .ZN(n_3066));
   NAND2_X1 i_2071 (.A1(in1[9]), .A2(in2[9]), .ZN(n_3067));
   OAI21_X1 i_2072 (.A(n_3065), .B1(n_3066), .B2(n_3067), .ZN(n_1626));
   NAND4_X1 i_2073 (.A1(in1[14]), .A2(in1[13]), .A3(in2[4]), .A4(in2[5]), 
      .ZN(n_3068));
   AOI22_X1 i_2074 (.A1(in1[14]), .A2(in2[4]), .B1(in1[13]), .B2(in2[5]), 
      .ZN(n_3070));
   NAND2_X1 i_2075 (.A1(in1[12]), .A2(in2[6]), .ZN(n_3071));
   OAI21_X1 i_2076 (.A(n_3068), .B1(n_3070), .B2(n_3071), .ZN(n_1633));
   INV_X1 i_2077 (.A(n_3047), .ZN(n_3072));
   NAND2_X1 i_2078 (.A1(n_3072), .A2(n_3051), .ZN(n_3073));
   XOR2_X1 i_2079 (.A(n_3073), .B(n_3048), .Z(n_1646));
   INV_X1 i_2080 (.A(n_3053), .ZN(n_3074));
   NAND2_X1 i_2081 (.A1(n_3074), .A2(n_3052), .ZN(n_3075));
   XOR2_X1 i_2082 (.A(n_3075), .B(n_3054), .Z(n_1604));
   INV_X1 i_2083 (.A(n_3058), .ZN(n_3114));
   NAND2_X1 i_2084 (.A1(n_3055), .A2(n_3114), .ZN(n_3117));
   XOR2_X1 i_2085 (.A(n_3117), .B(n_3059), .Z(n_1611));
   INV_X1 i_2086 (.A(n_3061), .ZN(n_3118));
   NAND2_X1 i_2087 (.A1(n_3118), .A2(n_3060), .ZN(n_3119));
   XOR2_X1 i_2088 (.A(n_3119), .B(n_3062), .Z(n_1618));
   INV_X1 i_2089 (.A(n_3066), .ZN(n_3120));
   NAND2_X1 i_2090 (.A1(n_3120), .A2(n_3065), .ZN(n_3121));
   XOR2_X1 i_2091 (.A(n_3121), .B(n_3067), .Z(n_1625));
   INV_X1 i_2092 (.A(n_3070), .ZN(n_3122));
   NAND2_X1 i_2093 (.A1(n_3122), .A2(n_3068), .ZN(n_3123));
   XOR2_X1 i_2094 (.A(n_3123), .B(n_3071), .Z(n_1632));
   INV_X1 i_2095 (.A(n_2944), .ZN(n_3126));
   NAND2_X1 i_2096 (.A1(n_3126), .A2(n_2943), .ZN(n_3127));
   XOR2_X1 i_2097 (.A(n_3127), .B(n_2945), .Z(n_1639));
   NAND4_X1 i_2098 (.A1(in2[16]), .A2(in2[15]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3128));
   AOI22_X1 i_2099 (.A1(in2[15]), .A2(in1[2]), .B1(in2[16]), .B2(in1[1]), 
      .ZN(n_3129));
   NAND2_X1 i_2100 (.A1(in2[17]), .A2(in1[0]), .ZN(n_3130));
   OAI21_X1 i_2101 (.A(n_3128), .B1(n_3129), .B2(n_3130), .ZN(n_1543));
   NOR2_X1 i_2102 (.A1(n_2262), .A2(n_598), .ZN(n_3133));
   NAND3_X1 i_2103 (.A1(n_3133), .A2(in2[13]), .A3(in1[4]), .ZN(n_3134));
   AOI21_X1 i_2104 (.A(n_3133), .B1(in2[13]), .B2(in1[4]), .ZN(n_3135));
   NAND2_X1 i_2105 (.A1(in2[14]), .A2(in1[3]), .ZN(n_3136));
   OAI21_X1 i_2106 (.A(n_3134), .B1(n_3135), .B2(n_3136), .ZN(n_1550));
   NAND4_X1 i_2107 (.A1(in2[10]), .A2(in1[8]), .A3(in2[9]), .A4(in1[7]), 
      .ZN(n_3137));
   AOI22_X1 i_2108 (.A1(in1[8]), .A2(in2[9]), .B1(in2[10]), .B2(in1[7]), 
      .ZN(n_3140));
   NAND2_X1 i_2109 (.A1(in2[11]), .A2(in1[6]), .ZN(n_3141));
   OAI21_X1 i_2110 (.A(n_3137), .B1(n_3140), .B2(n_3141), .ZN(n_1557));
   NAND4_X1 i_2111 (.A1(in1[11]), .A2(in1[10]), .A3(in2[7]), .A4(in2[6]), 
      .ZN(n_3142));
   AOI22_X1 i_2112 (.A1(in1[11]), .A2(in2[6]), .B1(in1[10]), .B2(in2[7]), 
      .ZN(n_3143));
   NAND2_X1 i_2113 (.A1(in1[9]), .A2(in2[8]), .ZN(n_3144));
   OAI21_X1 i_2114 (.A(n_3142), .B1(n_3143), .B2(n_3144), .ZN(n_1564));
   INV_X1 i_2115 (.A(n_3129), .ZN(n_3147));
   NAND2_X1 i_2116 (.A1(n_3147), .A2(n_3128), .ZN(n_3148));
   XOR2_X1 i_2117 (.A(n_3148), .B(n_3130), .Z(n_1542));
   INV_X1 i_2118 (.A(n_3135), .ZN(n_3149));
   NAND2_X1 i_2119 (.A1(n_3134), .A2(n_3149), .ZN(n_3150));
   XOR2_X1 i_2120 (.A(n_3150), .B(n_3136), .Z(n_1549));
   INV_X1 i_2121 (.A(n_3140), .ZN(n_3151));
   NAND2_X1 i_2122 (.A1(n_3151), .A2(n_3137), .ZN(n_3154));
   XOR2_X1 i_2123 (.A(n_3154), .B(n_3141), .Z(n_1556));
   INV_X1 i_2124 (.A(n_3143), .ZN(n_3155));
   NAND2_X1 i_2125 (.A1(n_3155), .A2(n_3142), .ZN(n_3156));
   XOR2_X1 i_2126 (.A(n_3156), .B(n_3144), .Z(n_1563));
   INV_X1 i_2127 (.A(n_3038), .ZN(n_3157));
   NAND2_X1 i_2128 (.A1(n_3157), .A2(n_3037), .ZN(n_3158));
   XOR2_X1 i_2129 (.A(n_3158), .B(n_3039), .Z(n_1570));
   INV_X1 i_2130 (.A(n_3044), .ZN(n_3161));
   NAND2_X1 i_2131 (.A1(n_3161), .A2(n_3041), .ZN(n_3162));
   XOR2_X1 i_2132 (.A(n_3162), .B(n_3045), .Z(n_1577));
   NAND4_X1 i_2133 (.A1(in1[14]), .A2(in1[13]), .A3(in2[2]), .A4(in2[1]), 
      .ZN(n_3163));
   AOI22_X1 i_2134 (.A1(in1[14]), .A2(in2[1]), .B1(in1[13]), .B2(in2[2]), 
      .ZN(n_3164));
   NAND2_X1 i_2135 (.A1(in1[12]), .A2(in2[3]), .ZN(n_3165));
   OAI21_X1 i_2136 (.A(n_3163), .B1(n_3164), .B2(n_3165), .ZN(n_3168));
   AOI21_X1 i_2137 (.A(n_3168), .B1(in1[16]), .B2(in2[0]), .ZN(n_3169));
   NAND2_X1 i_2138 (.A1(in1[15]), .A2(in2[1]), .ZN(n_3170));
   NAND3_X1 i_2139 (.A1(n_3168), .A2(in1[16]), .A3(in2[0]), .ZN(n_3171));
   AOI21_X1 i_2140 (.A(n_3169), .B1(n_3170), .B2(n_3171), .ZN(n_1516));
   NAND4_X1 i_2141 (.A1(in2[15]), .A2(in2[14]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3172));
   AOI22_X1 i_2142 (.A1(in2[14]), .A2(in1[2]), .B1(in2[15]), .B2(in1[1]), 
      .ZN(n_3175));
   NAND2_X1 i_2143 (.A1(in2[16]), .A2(in1[0]), .ZN(n_3176));
   OAI21_X1 i_2144 (.A(n_3172), .B1(n_3175), .B2(n_3176), .ZN(n_1482));
   NOR2_X1 i_2145 (.A1(n_2259), .A2(n_598), .ZN(n_3177));
   NAND3_X1 i_2146 (.A1(n_3177), .A2(in2[12]), .A3(in1[4]), .ZN(n_3178));
   AOI21_X1 i_2147 (.A(n_3177), .B1(in2[12]), .B2(in1[4]), .ZN(n_3179));
   NAND2_X1 i_2148 (.A1(in2[13]), .A2(in1[3]), .ZN(n_3182));
   OAI21_X1 i_2149 (.A(n_3178), .B1(n_3179), .B2(n_3182), .ZN(n_1489));
   NAND4_X1 i_2150 (.A1(in1[8]), .A2(in2[9]), .A3(in2[8]), .A4(in1[7]), .ZN(
      n_3183));
   AOI22_X1 i_2151 (.A1(in1[8]), .A2(in2[8]), .B1(in2[9]), .B2(in1[7]), .ZN(
      n_3184));
   NAND2_X1 i_2152 (.A1(in2[10]), .A2(in1[6]), .ZN(n_3185));
   OAI21_X1 i_2153 (.A(n_3183), .B1(n_3184), .B2(n_3185), .ZN(n_1496));
   NAND4_X1 i_2154 (.A1(in1[11]), .A2(in1[10]), .A3(in2[6]), .A4(in2[5]), 
      .ZN(n_3222));
   AOI22_X1 i_2155 (.A1(in1[11]), .A2(in2[5]), .B1(in1[10]), .B2(in2[6]), 
      .ZN(n_3225));
   NAND2_X1 i_2156 (.A1(in1[9]), .A2(in2[7]), .ZN(n_3226));
   OAI21_X1 i_2157 (.A(n_3222), .B1(n_3225), .B2(n_3226), .ZN(n_1503));
   NAND4_X1 i_2158 (.A1(in1[14]), .A2(in1[13]), .A3(in2[2]), .A4(in2[3]), 
      .ZN(n_3227));
   AOI22_X1 i_2159 (.A1(in1[14]), .A2(in2[2]), .B1(in1[13]), .B2(in2[3]), 
      .ZN(n_3228));
   NAND2_X1 i_2160 (.A1(in1[12]), .A2(in2[4]), .ZN(n_3229));
   OAI21_X1 i_2161 (.A(n_3227), .B1(n_3228), .B2(n_3229), .ZN(n_1510));
   INV_X1 i_2162 (.A(n_3175), .ZN(n_3230));
   NAND2_X1 i_2163 (.A1(n_3230), .A2(n_3172), .ZN(n_3231));
   XOR2_X1 i_2164 (.A(n_3231), .B(n_3176), .Z(n_1481));
   INV_X1 i_2165 (.A(n_3179), .ZN(n_3234));
   NAND2_X1 i_2166 (.A1(n_3178), .A2(n_3234), .ZN(n_3235));
   XOR2_X1 i_2167 (.A(n_3235), .B(n_3182), .Z(n_1488));
   INV_X1 i_2168 (.A(n_3184), .ZN(n_3236));
   NAND2_X1 i_2169 (.A1(n_3236), .A2(n_3183), .ZN(n_3237));
   XOR2_X1 i_2170 (.A(n_3237), .B(n_3185), .Z(n_1495));
   INV_X1 i_2171 (.A(n_3225), .ZN(n_3238));
   NAND2_X1 i_2172 (.A1(n_3238), .A2(n_3222), .ZN(n_3241));
   XOR2_X1 i_2173 (.A(n_3241), .B(n_3226), .Z(n_1502));
   INV_X1 i_2174 (.A(n_3228), .ZN(n_3242));
   NAND2_X1 i_2175 (.A1(n_3242), .A2(n_3227), .ZN(n_3243));
   XOR2_X1 i_2176 (.A(n_3243), .B(n_3229), .Z(n_1509));
   INV_X1 i_2177 (.A(n_3169), .ZN(n_3244));
   NAND2_X1 i_2178 (.A1(n_3244), .A2(n_3171), .ZN(n_3245));
   XOR2_X1 i_2179 (.A(n_3245), .B(n_3170), .Z(n_1515));
   NAND4_X1 i_2180 (.A1(in1[11]), .A2(in1[10]), .A3(in2[3]), .A4(in2[4]), 
      .ZN(n_3248));
   AOI22_X1 i_2181 (.A1(in1[11]), .A2(in2[3]), .B1(in1[10]), .B2(in2[4]), 
      .ZN(n_3249));
   NAND2_X1 i_2182 (.A1(in1[9]), .A2(in2[5]), .ZN(n_3250));
   OAI21_X1 i_2183 (.A(n_3248), .B1(n_3249), .B2(n_3250), .ZN(n_3251));
   NAND4_X1 i_2184 (.A1(in1[14]), .A2(in1[13]), .A3(in2[1]), .A4(in2[0]), 
      .ZN(n_3252));
   AOI22_X1 i_2185 (.A1(in1[14]), .A2(in2[0]), .B1(in1[13]), .B2(in2[1]), 
      .ZN(n_3255));
   NAND2_X1 i_2186 (.A1(in1[12]), .A2(in2[2]), .ZN(n_3256));
   OAI21_X1 i_2187 (.A(n_3252), .B1(n_3255), .B2(n_3256), .ZN(n_3257));
   NOR2_X1 i_2188 (.A1(n_3251), .A2(n_3257), .ZN(n_3258));
   NAND2_X1 i_2189 (.A1(in1[15]), .A2(in2[0]), .ZN(n_3259));
   NAND2_X1 i_2190 (.A1(n_3251), .A2(n_3257), .ZN(n_3262));
   AOI21_X1 i_2191 (.A(n_3258), .B1(n_3259), .B2(n_3262), .ZN(n_1458));
   NAND4_X1 i_2192 (.A1(in2[14]), .A2(in2[13]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3263));
   AOI22_X1 i_2193 (.A1(in2[13]), .A2(in1[2]), .B1(in2[14]), .B2(in1[1]), 
      .ZN(n_3264));
   NAND2_X1 i_2194 (.A1(in2[15]), .A2(in1[0]), .ZN(n_3265));
   OAI21_X1 i_2195 (.A(n_3263), .B1(n_3264), .B2(n_3265), .ZN(n_1423));
   NAND3_X1 i_2196 (.A1(n_3177), .A2(in2[10]), .A3(in1[4]), .ZN(n_3266));
   AOI22_X1 i_2197 (.A1(in2[10]), .A2(in1[5]), .B1(in2[11]), .B2(in1[4]), 
      .ZN(n_3269));
   NAND2_X1 i_2198 (.A1(in2[12]), .A2(in1[3]), .ZN(n_3270));
   OAI21_X1 i_2199 (.A(n_3266), .B1(n_3269), .B2(n_3270), .ZN(n_1430));
   NAND4_X1 i_2200 (.A1(in1[8]), .A2(in2[8]), .A3(in1[7]), .A4(in2[7]), .ZN(
      n_3271));
   AOI22_X1 i_2201 (.A1(in1[8]), .A2(in2[7]), .B1(in2[8]), .B2(in1[7]), .ZN(
      n_3272));
   NAND2_X1 i_2202 (.A1(in2[9]), .A2(in1[6]), .ZN(n_3273));
   OAI21_X1 i_2203 (.A(n_3271), .B1(n_3272), .B2(n_3273), .ZN(n_1437));
   NAND4_X1 i_2204 (.A1(in1[11]), .A2(in1[10]), .A3(in2[4]), .A4(in2[5]), 
      .ZN(n_3276));
   AOI22_X1 i_2205 (.A1(in1[11]), .A2(in2[4]), .B1(in1[10]), .B2(in2[5]), 
      .ZN(n_3277));
   NAND2_X1 i_2206 (.A1(in1[9]), .A2(in2[6]), .ZN(n_3278));
   OAI21_X1 i_2207 (.A(n_3276), .B1(n_3277), .B2(n_3278), .ZN(n_1444));
   INV_X1 i_2208 (.A(n_3258), .ZN(n_3279));
   NAND2_X1 i_2209 (.A1(n_3279), .A2(n_3262), .ZN(n_3280));
   XOR2_X1 i_2210 (.A(n_3280), .B(n_3259), .Z(n_1457));
   INV_X1 i_2211 (.A(n_3264), .ZN(n_3283));
   NAND2_X1 i_2212 (.A1(n_3283), .A2(n_3263), .ZN(n_3284));
   XOR2_X1 i_2213 (.A(n_3284), .B(n_3265), .Z(n_1422));
   INV_X1 i_2214 (.A(n_3269), .ZN(n_3285));
   NAND2_X1 i_2215 (.A1(n_3266), .A2(n_3285), .ZN(n_3322));
   XOR2_X1 i_2216 (.A(n_3322), .B(n_3270), .Z(n_1429));
   INV_X1 i_2217 (.A(n_3272), .ZN(n_3325));
   NAND2_X1 i_2218 (.A1(n_3325), .A2(n_3271), .ZN(n_3326));
   XOR2_X1 i_2219 (.A(n_3326), .B(n_3273), .Z(n_1436));
   INV_X1 i_2220 (.A(n_3277), .ZN(n_3327));
   NAND2_X1 i_2221 (.A1(n_3327), .A2(n_3276), .ZN(n_3328));
   XOR2_X1 i_2222 (.A(n_3328), .B(n_3278), .Z(n_1443));
   INV_X1 i_2223 (.A(n_3164), .ZN(n_3329));
   NAND2_X1 i_2224 (.A1(n_3329), .A2(n_3163), .ZN(n_3330));
   XOR2_X1 i_2225 (.A(n_3330), .B(n_3165), .Z(n_1450));
   NAND4_X1 i_2226 (.A1(in2[13]), .A2(in2[12]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3331));
   AOI22_X1 i_2227 (.A1(in2[12]), .A2(in1[2]), .B1(in2[13]), .B2(in1[1]), 
      .ZN(n_3334));
   NAND2_X1 i_2228 (.A1(in2[14]), .A2(in1[0]), .ZN(n_3335));
   OAI21_X1 i_2229 (.A(n_3331), .B1(n_3334), .B2(n_3335), .ZN(n_1372));
   NOR2_X1 i_2230 (.A1(n_996), .A2(n_598), .ZN(n_3336));
   NAND3_X1 i_2231 (.A1(n_3336), .A2(in2[10]), .A3(in1[4]), .ZN(n_3337));
   AOI21_X1 i_2232 (.A(n_3336), .B1(in2[10]), .B2(in1[4]), .ZN(n_3338));
   NAND2_X1 i_2233 (.A1(in2[11]), .A2(in1[3]), .ZN(n_3341));
   OAI21_X1 i_2234 (.A(n_3337), .B1(n_3338), .B2(n_3341), .ZN(n_1379));
   NAND4_X1 i_2235 (.A1(in1[8]), .A2(in1[7]), .A3(in2[7]), .A4(in2[6]), .ZN(
      n_3342));
   AOI22_X1 i_2236 (.A1(in1[8]), .A2(in2[6]), .B1(in1[7]), .B2(in2[7]), .ZN(
      n_3343));
   NAND2_X1 i_2237 (.A1(in2[8]), .A2(in1[6]), .ZN(n_3344));
   OAI21_X1 i_2238 (.A(n_3342), .B1(n_3343), .B2(n_3344), .ZN(n_1386));
   INV_X1 i_2239 (.A(n_3334), .ZN(n_3345));
   NAND2_X1 i_2240 (.A1(n_3345), .A2(n_3331), .ZN(n_3348));
   XOR2_X1 i_2241 (.A(n_3348), .B(n_3335), .Z(n_1371));
   INV_X1 i_2242 (.A(n_3338), .ZN(n_3349));
   NAND2_X1 i_2243 (.A1(n_3337), .A2(n_3349), .ZN(n_3350));
   XOR2_X1 i_2244 (.A(n_3350), .B(n_3341), .Z(n_1378));
   INV_X1 i_2245 (.A(n_3343), .ZN(n_3351));
   NAND2_X1 i_2246 (.A1(n_3351), .A2(n_3342), .ZN(n_3352));
   XOR2_X1 i_2247 (.A(n_3352), .B(n_3344), .Z(n_1385));
   INV_X1 i_2248 (.A(n_3249), .ZN(n_3355));
   NAND2_X1 i_2249 (.A1(n_3355), .A2(n_3248), .ZN(n_3356));
   XOR2_X1 i_2250 (.A(n_3356), .B(n_3250), .Z(n_1392));
   INV_X1 i_2251 (.A(n_3255), .ZN(n_3357));
   NAND2_X1 i_2252 (.A1(n_3357), .A2(n_3252), .ZN(n_3358));
   XOR2_X1 i_2253 (.A(n_3358), .B(n_3256), .Z(n_1399));
   NAND4_X1 i_2254 (.A1(in1[11]), .A2(in1[10]), .A3(in2[2]), .A4(in2[1]), 
      .ZN(n_3359));
   AOI22_X1 i_2255 (.A1(in1[11]), .A2(in2[1]), .B1(in1[10]), .B2(in2[2]), 
      .ZN(n_3362));
   NAND2_X1 i_2256 (.A1(in1[9]), .A2(in2[3]), .ZN(n_3363));
   OAI21_X1 i_2257 (.A(n_3359), .B1(n_3362), .B2(n_3363), .ZN(n_3364));
   AOI21_X1 i_2258 (.A(n_3364), .B1(in1[13]), .B2(in2[0]), .ZN(n_3365));
   NAND2_X1 i_2259 (.A1(in1[12]), .A2(in2[1]), .ZN(n_3366));
   NAND3_X1 i_2260 (.A1(n_3364), .A2(in1[13]), .A3(in2[0]), .ZN(n_3369));
   AOI21_X1 i_2261 (.A(n_3365), .B1(n_3366), .B2(n_3369), .ZN(n_1349));
   NAND4_X1 i_2262 (.A1(in2[12]), .A2(in2[11]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3370));
   AOI22_X1 i_2263 (.A1(in2[11]), .A2(in1[2]), .B1(in2[12]), .B2(in1[1]), 
      .ZN(n_3371));
   NAND2_X1 i_2264 (.A1(in2[13]), .A2(in1[0]), .ZN(n_3372));
   OAI21_X1 i_2265 (.A(n_3370), .B1(n_3371), .B2(n_3372), .ZN(n_1322));
   NOR2_X1 i_2266 (.A1(n_994), .A2(n_598), .ZN(n_3373));
   NAND3_X1 i_2267 (.A1(n_3373), .A2(in2[9]), .A3(in1[4]), .ZN(n_3376));
   AOI21_X1 i_2268 (.A(n_3373), .B1(in2[9]), .B2(in1[4]), .ZN(n_3377));
   NAND2_X1 i_2269 (.A1(in2[10]), .A2(in1[3]), .ZN(n_3378));
   OAI21_X1 i_2270 (.A(n_3376), .B1(n_3377), .B2(n_3378), .ZN(n_1329));
   NAND4_X1 i_2271 (.A1(in1[8]), .A2(in1[7]), .A3(in2[6]), .A4(in2[5]), .ZN(
      n_3379));
   AOI22_X1 i_2272 (.A1(in1[8]), .A2(in2[5]), .B1(in1[7]), .B2(in2[6]), .ZN(
      n_3381));
   NAND2_X1 i_2273 (.A1(in2[7]), .A2(in1[6]), .ZN(n_3382));
   OAI21_X1 i_2274 (.A(n_3379), .B1(n_3381), .B2(n_3382), .ZN(n_1336));
   NAND4_X1 i_2275 (.A1(in1[11]), .A2(in1[10]), .A3(in2[2]), .A4(in2[3]), 
      .ZN(n_3383));
   AOI22_X1 i_2276 (.A1(in1[11]), .A2(in2[2]), .B1(in1[10]), .B2(in2[3]), 
      .ZN(n_3384));
   NAND2_X1 i_2277 (.A1(in1[9]), .A2(in2[4]), .ZN(n_3385));
   OAI21_X1 i_2278 (.A(n_3383), .B1(n_3384), .B2(n_3385), .ZN(n_1343));
   INV_X1 i_2279 (.A(n_3371), .ZN(n_3386));
   NAND2_X1 i_2280 (.A1(n_3386), .A2(n_3370), .ZN(n_3421));
   XOR2_X1 i_2281 (.A(n_3421), .B(n_3372), .Z(n_1321));
   INV_X1 i_2282 (.A(n_3377), .ZN(n_3424));
   NAND2_X1 i_2283 (.A1(n_3376), .A2(n_3424), .ZN(n_3425));
   XOR2_X1 i_2284 (.A(n_3425), .B(n_3378), .Z(n_1328));
   INV_X1 i_2285 (.A(n_3381), .ZN(n_3426));
   NAND2_X1 i_2286 (.A1(n_3426), .A2(n_3379), .ZN(n_3427));
   XOR2_X1 i_2287 (.A(n_3427), .B(n_3382), .Z(n_1335));
   INV_X1 i_2288 (.A(n_3384), .ZN(n_3428));
   NAND2_X1 i_2289 (.A1(n_3428), .A2(n_3383), .ZN(n_3429));
   XOR2_X1 i_2290 (.A(n_3429), .B(n_3385), .Z(n_1342));
   INV_X1 i_2291 (.A(n_3365), .ZN(n_3430));
   NAND2_X1 i_2292 (.A1(n_3430), .A2(n_3369), .ZN(n_3433));
   XOR2_X1 i_2293 (.A(n_3433), .B(n_3366), .Z(n_1348));
   NAND4_X1 i_2294 (.A1(in1[8]), .A2(in1[7]), .A3(in2[3]), .A4(in2[4]), .ZN(
      n_3434));
   AOI22_X1 i_2295 (.A1(in1[8]), .A2(in2[3]), .B1(in1[7]), .B2(in2[4]), .ZN(
      n_3435));
   NAND2_X1 i_2296 (.A1(in1[6]), .A2(in2[5]), .ZN(n_3436));
   OAI21_X1 i_2297 (.A(n_3434), .B1(n_3435), .B2(n_3436), .ZN(n_3437));
   NAND4_X1 i_2298 (.A1(in1[11]), .A2(in1[10]), .A3(in2[1]), .A4(in2[0]), 
      .ZN(n_3440));
   AOI22_X1 i_2299 (.A1(in1[11]), .A2(in2[0]), .B1(in1[10]), .B2(in2[1]), 
      .ZN(n_3441));
   NAND2_X1 i_2300 (.A1(in1[9]), .A2(in2[2]), .ZN(n_3442));
   OAI21_X1 i_2301 (.A(n_3440), .B1(n_3441), .B2(n_3442), .ZN(n_3443));
   NOR2_X1 i_2302 (.A1(n_3437), .A2(n_3443), .ZN(n_3444));
   NAND2_X1 i_2303 (.A1(in1[12]), .A2(in2[0]), .ZN(n_3447));
   NAND2_X1 i_2304 (.A1(n_3437), .A2(n_3443), .ZN(n_3448));
   AOI21_X1 i_2305 (.A(n_3444), .B1(n_3447), .B2(n_3448), .ZN(n_1302));
   NAND4_X1 i_2306 (.A1(in2[11]), .A2(in2[10]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3449));
   AOI22_X1 i_2307 (.A1(in2[10]), .A2(in1[2]), .B1(in2[11]), .B2(in1[1]), 
      .ZN(n_3450));
   NAND2_X1 i_2308 (.A1(in2[12]), .A2(in1[0]), .ZN(n_3451));
   OAI21_X1 i_2309 (.A(n_3449), .B1(n_3450), .B2(n_3451), .ZN(n_1274));
   NAND3_X1 i_2310 (.A1(n_3373), .A2(in2[7]), .A3(in1[4]), .ZN(n_3454));
   AOI22_X1 i_2311 (.A1(in2[7]), .A2(in1[5]), .B1(in2[8]), .B2(in1[4]), .ZN(
      n_3455));
   NAND2_X1 i_2312 (.A1(in2[9]), .A2(in1[3]), .ZN(n_3456));
   OAI21_X1 i_2313 (.A(n_3454), .B1(n_3455), .B2(n_3456), .ZN(n_1281));
   NAND4_X1 i_2314 (.A1(in1[8]), .A2(in1[7]), .A3(in2[4]), .A4(in2[5]), .ZN(
      n_3457));
   AOI22_X1 i_2315 (.A1(in1[8]), .A2(in2[4]), .B1(in1[7]), .B2(in2[5]), .ZN(
      n_3458));
   NAND2_X1 i_2316 (.A1(in1[6]), .A2(in2[6]), .ZN(n_3461));
   OAI21_X1 i_2317 (.A(n_3457), .B1(n_3458), .B2(n_3461), .ZN(n_1288));
   INV_X1 i_2318 (.A(n_3444), .ZN(n_3462));
   NAND2_X1 i_2319 (.A1(n_3462), .A2(n_3448), .ZN(n_3463));
   XOR2_X1 i_2320 (.A(n_3463), .B(n_3447), .Z(n_1301));
   INV_X1 i_2321 (.A(n_3450), .ZN(n_3464));
   NAND2_X1 i_2322 (.A1(n_3464), .A2(n_3449), .ZN(n_3465));
   XOR2_X1 i_2323 (.A(n_3465), .B(n_3451), .Z(n_1273));
   INV_X1 i_2324 (.A(n_3455), .ZN(n_3468));
   NAND2_X1 i_2325 (.A1(n_3454), .A2(n_3468), .ZN(n_3469));
   XOR2_X1 i_2326 (.A(n_3469), .B(n_3456), .Z(n_1280));
   INV_X1 i_2327 (.A(n_3458), .ZN(n_3470));
   NAND2_X1 i_2328 (.A1(n_3470), .A2(n_3457), .ZN(n_3471));
   XOR2_X1 i_2329 (.A(n_3471), .B(n_3461), .Z(n_1287));
   INV_X1 i_2330 (.A(n_3362), .ZN(n_3472));
   NAND2_X1 i_2331 (.A1(n_3472), .A2(n_3359), .ZN(n_3475));
   XOR2_X1 i_2332 (.A(n_3475), .B(n_3363), .Z(n_1294));
   NAND4_X1 i_2333 (.A1(in2[10]), .A2(in2[9]), .A3(in1[2]), .A4(in1[1]), 
      .ZN(n_3476));
   AOI22_X1 i_2334 (.A1(in2[9]), .A2(in1[2]), .B1(in2[10]), .B2(in1[1]), 
      .ZN(n_3477));
   NAND2_X1 i_2335 (.A1(in2[11]), .A2(in1[0]), .ZN(n_3478));
   OAI21_X1 i_2336 (.A(n_3476), .B1(n_3477), .B2(n_3478), .ZN(n_1234));
   NOR2_X1 i_2337 (.A1(n_598), .A2(n_2083), .ZN(n_3479));
   NAND3_X1 i_2338 (.A1(n_3479), .A2(in2[7]), .A3(in1[4]), .ZN(n_3482));
   AOI21_X1 i_2339 (.A(n_3479), .B1(in2[7]), .B2(in1[4]), .ZN(n_3483));
   NAND2_X1 i_2340 (.A1(in2[8]), .A2(in1[3]), .ZN(n_3484));
   OAI21_X1 i_2341 (.A(n_3482), .B1(n_3483), .B2(n_3484), .ZN(n_1241));
   INV_X1 i_2342 (.A(n_3477), .ZN(n_3485));
   NAND2_X1 i_2343 (.A1(n_3485), .A2(n_3476), .ZN(n_3518));
   XOR2_X1 i_2344 (.A(n_3518), .B(n_3478), .Z(n_1233));
   INV_X1 i_2345 (.A(n_3483), .ZN(n_3521));
   NAND2_X1 i_2346 (.A1(n_3482), .A2(n_3521), .ZN(n_3522));
   XOR2_X1 i_2347 (.A(n_3522), .B(n_3484), .Z(n_1240));
   INV_X1 i_2348 (.A(n_3435), .ZN(n_3523));
   NAND2_X1 i_2349 (.A1(n_3523), .A2(n_3434), .ZN(n_3524));
   XOR2_X1 i_2350 (.A(n_3524), .B(n_3436), .Z(n_1247));
   INV_X1 i_2351 (.A(n_3441), .ZN(n_3525));
   NAND2_X1 i_2352 (.A1(n_3525), .A2(n_3440), .ZN(n_3526));
   XOR2_X1 i_2353 (.A(n_3526), .B(n_3442), .Z(n_1254));
   NAND4_X1 i_2354 (.A1(in1[8]), .A2(in2[2]), .A3(in1[7]), .A4(in2[1]), .ZN(
      n_3527));
   AOI22_X1 i_2355 (.A1(in1[8]), .A2(in2[1]), .B1(in2[2]), .B2(in1[7]), .ZN(
      n_3530));
   NAND2_X1 i_2356 (.A1(in2[3]), .A2(in1[6]), .ZN(n_3531));
   OAI21_X1 i_2357 (.A(n_3527), .B1(n_3530), .B2(n_3531), .ZN(n_3532));
   AOI21_X1 i_2358 (.A(n_3532), .B1(in1[10]), .B2(in2[0]), .ZN(n_3533));
   NAND2_X1 i_2359 (.A1(in1[9]), .A2(in2[1]), .ZN(n_3534));
   NAND3_X1 i_2360 (.A1(n_3532), .A2(in1[10]), .A3(in2[0]), .ZN(n_3537));
   AOI21_X1 i_2361 (.A(n_3533), .B1(n_3534), .B2(n_3537), .ZN(n_1215));
   NAND4_X1 i_2362 (.A1(in2[9]), .A2(in2[8]), .A3(in1[2]), .A4(in1[1]), .ZN(
      n_3538));
   AOI22_X1 i_2363 (.A1(in2[8]), .A2(in1[2]), .B1(in2[9]), .B2(in1[1]), .ZN(
      n_3539));
   NAND2_X1 i_2364 (.A1(in2[10]), .A2(in1[0]), .ZN(n_3540));
   OAI21_X1 i_2365 (.A(n_3538), .B1(n_3539), .B2(n_3540), .ZN(n_1195));
   NOR2_X1 i_2366 (.A1(n_598), .A2(n_694), .ZN(n_3541));
   NAND3_X1 i_2367 (.A1(n_3541), .A2(in1[4]), .A3(in2[6]), .ZN(n_3544));
   AOI21_X1 i_2368 (.A(n_3541), .B1(in1[4]), .B2(in2[6]), .ZN(n_3545));
   NAND2_X1 i_2369 (.A1(in2[7]), .A2(in1[3]), .ZN(n_3546));
   OAI21_X1 i_2370 (.A(n_3544), .B1(n_3545), .B2(n_3546), .ZN(n_1202));
   NAND4_X1 i_2371 (.A1(in1[8]), .A2(in2[2]), .A3(in1[7]), .A4(in2[3]), .ZN(
      n_3547));
   AOI22_X1 i_2372 (.A1(in1[8]), .A2(in2[2]), .B1(in1[7]), .B2(in2[3]), .ZN(
      n_3548));
   NAND2_X1 i_2373 (.A1(in1[6]), .A2(in2[4]), .ZN(n_3551));
   OAI21_X1 i_2374 (.A(n_3547), .B1(n_3548), .B2(n_3551), .ZN(n_1209));
   INV_X1 i_2375 (.A(n_3539), .ZN(n_3552));
   NAND2_X1 i_2376 (.A1(n_3552), .A2(n_3538), .ZN(n_3553));
   XOR2_X1 i_2377 (.A(n_3553), .B(n_3540), .Z(n_1194));
   INV_X1 i_2378 (.A(n_3545), .ZN(n_3554));
   NAND2_X1 i_2379 (.A1(n_3544), .A2(n_3554), .ZN(n_3555));
   XOR2_X1 i_2380 (.A(n_3555), .B(n_3546), .Z(n_1201));
   INV_X1 i_2381 (.A(n_3548), .ZN(n_3558));
   NAND2_X1 i_2382 (.A1(n_3558), .A2(n_3547), .ZN(n_3559));
   XOR2_X1 i_2383 (.A(n_3559), .B(n_3551), .Z(n_1208));
   INV_X1 i_2384 (.A(n_3533), .ZN(n_3560));
   NAND2_X1 i_2385 (.A1(n_3560), .A2(n_3537), .ZN(n_3561));
   XOR2_X1 i_2386 (.A(n_3561), .B(n_3534), .Z(n_1214));
   AOI21_X1 i_2387 (.A(n_575), .B1(n_574), .B2(n_576), .ZN(n_1179));
   NAND4_X1 i_2388 (.A1(in2[8]), .A2(in2[7]), .A3(in1[2]), .A4(in1[1]), .ZN(
      n_3612));
   AOI22_X1 i_2389 (.A1(in2[7]), .A2(in1[2]), .B1(in2[8]), .B2(in1[1]), .ZN(
      n_3613));
   NAND2_X1 i_2390 (.A1(in2[9]), .A2(in1[0]), .ZN(n_3614));
   OAI21_X1 i_2391 (.A(n_3612), .B1(n_3613), .B2(n_3614), .ZN(n_1158));
   NAND3_X1 i_2392 (.A1(n_3541), .A2(in1[4]), .A3(in2[4]), .ZN(n_3615));
   AOI22_X1 i_2393 (.A1(in1[5]), .A2(in2[4]), .B1(in1[4]), .B2(in2[5]), .ZN(
      n_3616));
   NAND2_X1 i_2394 (.A1(in2[6]), .A2(in1[3]), .ZN(n_3619));
   OAI21_X1 i_2395 (.A(n_3615), .B1(n_3616), .B2(n_3619), .ZN(n_1165));
   INV_X1 i_2396 (.A(n_3613), .ZN(n_3622));
   NAND2_X1 i_2397 (.A1(n_3622), .A2(n_3612), .ZN(n_3623));
   XOR2_X1 i_2398 (.A(n_3623), .B(n_3614), .Z(n_1157));
   INV_X1 i_2399 (.A(n_3616), .ZN(n_3626));
   NAND2_X1 i_2400 (.A1(n_3615), .A2(n_3626), .ZN(n_3627));
   XOR2_X1 i_2401 (.A(n_3627), .B(n_3619), .Z(n_1164));
   INV_X1 i_2402 (.A(n_3530), .ZN(n_3628));
   NAND2_X1 i_2403 (.A1(n_3628), .A2(n_3527), .ZN(n_3629));
   XOR2_X1 i_2404 (.A(n_3629), .B(n_3531), .Z(n_1171));
   NAND4_X1 i_2405 (.A1(in2[7]), .A2(in2[6]), .A3(in1[2]), .A4(in1[1]), .ZN(
      n_3630));
   AOI22_X1 i_2406 (.A1(in2[6]), .A2(in1[2]), .B1(in2[7]), .B2(in1[1]), .ZN(
      n_3633));
   NAND2_X1 i_2407 (.A1(in2[8]), .A2(in1[0]), .ZN(n_3634));
   OAI21_X1 i_2408 (.A(n_3630), .B1(n_3633), .B2(n_3634), .ZN(n_1129));
   INV_X1 i_2409 (.A(n_3633), .ZN(n_3635));
   NAND2_X1 i_2410 (.A1(n_3635), .A2(n_3630), .ZN(n_3636));
   XOR2_X1 i_2411 (.A(n_3636), .B(n_3634), .Z(n_1128));
   INV_X1 i_2412 (.A(n_596), .ZN(n_3637));
   NAND2_X1 i_2413 (.A1(n_597), .A2(n_3637), .ZN(n_3640));
   XOR2_X1 i_2414 (.A(n_3640), .B(n_595), .Z(n_1135));
   INV_X1 i_2415 (.A(n_593), .ZN(n_3641));
   NAND2_X1 i_2416 (.A1(n_3641), .A2(n_594), .ZN(n_3642));
   XOR2_X1 i_2417 (.A(n_3642), .B(n_579), .Z(n_1142));
   AOI21_X1 i_2418 (.A(n_659), .B1(n_656), .B2(n_658), .ZN(n_1114));
   NAND4_X1 i_2419 (.A1(in2[6]), .A2(in1[2]), .A3(in2[5]), .A4(in1[1]), .ZN(
      n_3657));
   AOI22_X1 i_2420 (.A1(in1[2]), .A2(in2[5]), .B1(in2[6]), .B2(in1[1]), .ZN(
      n_3659));
   NAND2_X1 i_2421 (.A1(in2[7]), .A2(in1[0]), .ZN(n_3660));
   OAI21_X1 i_2422 (.A(n_3657), .B1(n_3659), .B2(n_3660), .ZN(n_1101));
   INV_X1 i_2423 (.A(n_664), .ZN(n_3661));
   NAND3_X1 i_2424 (.A1(n_3661), .A2(in2[3]), .A3(in1[4]), .ZN(n_3662));
   AOI21_X1 i_2425 (.A(n_3661), .B1(in2[3]), .B2(in1[4]), .ZN(n_3663));
   NAND2_X1 i_2426 (.A1(in2[4]), .A2(in1[3]), .ZN(n_3664));
   OAI21_X1 i_2427 (.A(n_3662), .B1(n_3663), .B2(n_3664), .ZN(n_1108));
   INV_X1 i_2428 (.A(n_3659), .ZN(n_3695));
   NAND2_X1 i_2429 (.A1(n_3695), .A2(n_3657), .ZN(n_3698));
   XOR2_X1 i_2430 (.A(n_3698), .B(n_3660), .Z(n_1100));
   INV_X1 i_2431 (.A(n_3663), .ZN(n_3699));
   NAND2_X1 i_2432 (.A1(n_3662), .A2(n_3699), .ZN(n_3700));
   XOR2_X1 i_2433 (.A(n_3700), .B(n_3664), .Z(n_1107));
   NAND2_X1 i_2434 (.A1(n_677), .A2(n_675), .ZN(n_3735));
   XNOR2_X1 i_2435 (.A(n_3735), .B(n_676), .ZN(n_1056));
   NAND2_X1 i_2436 (.A1(n_672), .A2(n_669), .ZN(n_3736));
   XNOR2_X1 i_2437 (.A(n_3736), .B(n_670), .ZN(n_1063));
   INV_X1 i_2438 (.A(n_520), .ZN(n_3737));
   AOI21_X1 i_2439 (.A(n_521), .B1(n_3737), .B2(n_523), .ZN(n_1040));
   OAI21_X1 i_2440 (.A(n_539), .B1(n_527), .B2(n_673), .ZN(n_3738));
   NAND3_X1 i_2441 (.A1(n_3738), .A2(in1[3]), .A3(in2[1]), .ZN(n_404));
   AOI22_X1 i_2442 (.A1(n_3738), .A2(in2[0]), .B1(n_527), .B2(n_539), .ZN(n_405));
   OAI21_X1 i_2443 (.A(n_404), .B1(n_405), .B2(n_1857), .ZN(n_1045));
   INV_X1 i_2444 (.A(n_3738), .ZN(n_1046));
   OAI21_X1 i_2445 (.A(n_534), .B1(n_535), .B2(n_538), .ZN(n_1030));
   INV_X1 i_2446 (.A(n_531), .ZN(n_406));
   AOI22_X1 i_2447 (.A1(in2[1]), .A2(in1[0]), .B1(in2[0]), .B2(in1[1]), .ZN(
      n_411));
   NOR2_X1 i_2448 (.A1(n_406), .A2(n_411), .ZN(out[1]));
   INV_X1 i_2449 (.A(n_530), .ZN(n_475));
   NAND2_X1 i_2450 (.A1(n_475), .A2(n_532), .ZN(n_517));
   XOR2_X1 i_2451 (.A(n_517), .B(n_531), .Z(out[2]));
   INV_X1 i_2452 (.A(n_364), .ZN(n_519));
   INV_X1 i_2453 (.A(n_305), .ZN(n_524));
   OAI22_X1 i_2454 (.A1(n_519), .A2(n_305), .B1(n_524), .B2(n_364), .ZN(n_525));
   NOR2_X1 i_2455 (.A1(n_1384), .A2(n_1602), .ZN(n_526));
   XOR2_X1 i_2456 (.A(n_525), .B(n_526), .Z(out[62]));
   NAND2_X1 i_2457 (.A1(n_524), .A2(n_519), .ZN(n_540));
   AOI22_X1 i_2458 (.A1(n_540), .A2(n_526), .B1(n_305), .B2(n_364), .ZN(out[63]));
   XOR2_X1 i_2459 (.A(n_574), .B(n_573), .Z(n_572));
   OAI21_X1 i_2460 (.A(n_576), .B1(n_578), .B2(n_577), .ZN(n_573));
   NAND2_X1 i_2461 (.A1(in2[0]), .A2(in1[9]), .ZN(n_574));
   NOR2_X1 i_2462 (.A1(n_578), .A2(n_577), .ZN(n_575));
   NAND2_X1 i_2463 (.A1(n_578), .A2(n_577), .ZN(n_576));
   OAI21_X1 i_2464 (.A(n_594), .B1(n_593), .B2(n_579), .ZN(n_577));
   OAI21_X1 i_2465 (.A(n_597), .B1(n_596), .B2(n_595), .ZN(n_578));
   NAND2_X1 i_2466 (.A1(in2[2]), .A2(in1[6]), .ZN(n_579));
   AOI22_X1 i_2467 (.A1(in2[0]), .A2(in1[8]), .B1(in2[1]), .B2(in1[7]), .ZN(
      n_593));
   NAND4_X1 i_2468 (.A1(in2[0]), .A2(in1[8]), .A3(in2[1]), .A4(in1[7]), .ZN(
      n_594));
   NAND2_X1 i_2469 (.A1(in2[5]), .A2(in1[3]), .ZN(n_595));
   AOI22_X1 i_2470 (.A1(in2[3]), .A2(in1[5]), .B1(in2[4]), .B2(in1[4]), .ZN(
      n_596));
   NAND4_X1 i_2471 (.A1(in2[3]), .A2(in1[5]), .A3(in2[4]), .A4(in1[4]), .ZN(
      n_597));
   INV_X1 i_2472 (.A(in1[5]), .ZN(n_598));
   INV_X1 i_2473 (.A(in2[3]), .ZN(n_599));
   FA_X1 i_2474 (.A(n_1075), .B(n_1089), .CI(n_1113), .CO(n_600), .S(n_1120));
   FA_X1 i_2475 (.A(n_1081), .B(n_1074), .CI(n_1088), .CO(n_1095), .S(n_601));
   HA_X1 i_2476 (.A(n_1120), .B(n_1095), .CO(n_603), .S(n_602));
   XOR2_X1 i_2477 (.A(n_646), .B(n_604), .Z(n_1088));
   OAI21_X1 i_2478 (.A(n_648), .B1(n_650), .B2(n_649), .ZN(n_604));
   XOR2_X1 i_2479 (.A(n_651), .B(n_643), .Z(n_1074));
   OAI21_X1 i_2480 (.A(n_653), .B1(n_655), .B2(n_654), .ZN(n_643));
   XOR2_X1 i_2481 (.A(n_661), .B(n_644), .Z(n_1081));
   OAI21_X1 i_2482 (.A(n_662), .B1(n_674), .B2(n_664), .ZN(n_644));
   XNOR2_X1 i_2483 (.A(n_656), .B(n_645), .ZN(n_1113));
   NOR2_X1 i_2484 (.A1(n_659), .A2(n_657), .ZN(n_645));
   OAI22_X1 i_2485 (.A1(n_650), .A2(n_649), .B1(n_647), .B2(n_646), .ZN(n_1089));
   NAND2_X1 i_2486 (.A1(in2[0]), .A2(in1[6]), .ZN(n_646));
   INV_X1 i_2487 (.A(n_648), .ZN(n_647));
   NAND2_X1 i_2488 (.A1(n_650), .A2(n_649), .ZN(n_648));
   AOI21_X1 i_2489 (.A(n_678), .B1(n_676), .B2(n_675), .ZN(n_649));
   OAI21_X1 i_2490 (.A(n_669), .B1(n_671), .B2(n_670), .ZN(n_650));
   OAI21_X1 i_2491 (.A(n_653), .B1(n_652), .B2(n_651), .ZN(n_1075));
   NAND2_X1 i_2492 (.A1(in2[6]), .A2(in1[0]), .ZN(n_651));
   NOR2_X1 i_2493 (.A1(n_655), .A2(n_654), .ZN(n_652));
   NAND2_X1 i_2494 (.A1(n_655), .A2(n_654), .ZN(n_653));
   NOR2_X1 i_2495 (.A1(n_694), .A2(n_691), .ZN(n_654));
   AND2_X1 i_2496 (.A1(in2[4]), .A2(in1[2]), .ZN(n_655));
   NAND2_X1 i_2497 (.A1(in2[1]), .A2(in1[6]), .ZN(n_656));
   INV_X1 i_2498 (.A(n_658), .ZN(n_657));
   NAND3_X1 i_2499 (.A1(in2[0]), .A2(in1[7]), .A3(n_660), .ZN(n_658));
   AOI21_X1 i_2500 (.A(n_660), .B1(in2[0]), .B2(in1[7]), .ZN(n_659));
   OAI22_X1 i_2501 (.A1(n_674), .A2(n_664), .B1(n_663), .B2(n_661), .ZN(n_660));
   NAND2_X1 i_2502 (.A1(in2[3]), .A2(in1[3]), .ZN(n_661));
   INV_X1 i_2503 (.A(n_663), .ZN(n_662));
   AOI22_X1 i_2504 (.A1(in2[1]), .A2(in1[5]), .B1(in2[2]), .B2(in1[4]), .ZN(
      n_663));
   NAND2_X1 i_2505 (.A1(in2[2]), .A2(in1[5]), .ZN(n_664));
   OAI21_X1 i_2506 (.A(n_674), .B1(n_692), .B2(n_598), .ZN(n_669));
   AND2_X1 i_2507 (.A1(in2[2]), .A2(in1[3]), .ZN(n_670));
   INV_X1 i_2508 (.A(n_672), .ZN(n_671));
   NAND3_X1 i_2509 (.A1(in1[5]), .A2(n_673), .A3(in2[0]), .ZN(n_672));
   INV_X1 i_2510 (.A(n_674), .ZN(n_673));
   NAND2_X1 i_2511 (.A1(in2[1]), .A2(in1[4]), .ZN(n_674));
   OAI21_X1 i_2512 (.A(n_679), .B1(n_693), .B2(n_691), .ZN(n_675));
   NOR2_X1 i_2513 (.A1(n_694), .A2(n_690), .ZN(n_676));
   INV_X1 i_2514 (.A(n_678), .ZN(n_677));
   NOR3_X1 i_2515 (.A1(n_693), .A2(n_691), .A3(n_679), .ZN(n_678));
   NAND2_X1 i_2516 (.A1(in2[3]), .A2(in1[2]), .ZN(n_679));
   INV_X1 i_2517 (.A(in1[0]), .ZN(n_690));
   INV_X1 i_2518 (.A(in1[1]), .ZN(n_691));
   INV_X1 i_2519 (.A(in2[0]), .ZN(n_692));
   INV_X1 i_2520 (.A(in2[4]), .ZN(n_693));
   INV_X1 i_2521 (.A(in2[5]), .ZN(n_694));
   OAI21_X1 i_2522 (.A(n_696), .B1(n_707), .B2(n_698), .ZN(n_695));
   NAND2_X1 i_2523 (.A1(n_707), .A2(n_698), .ZN(n_696));
   NOR2_X1 i_2524 (.A1(n_707), .A2(n_698), .ZN(n_697));
   OAI21_X1 i_2525 (.A(n_710), .B1(n_709), .B2(n_708), .ZN(n_698));
   OAI21_X1 i_2526 (.A(n_713), .B1(n_712), .B2(n_711), .ZN(n_707));
   NAND2_X1 i_2527 (.A1(in1[24]), .A2(in2[2]), .ZN(n_708));
   AOI22_X1 i_2528 (.A1(in1[25]), .A2(in2[1]), .B1(in1[26]), .B2(in2[0]), 
      .ZN(n_709));
   NAND4_X1 i_2529 (.A1(in1[25]), .A2(in2[1]), .A3(in1[26]), .A4(in2[0]), 
      .ZN(n_710));
   NAND2_X1 i_2530 (.A1(in1[21]), .A2(in2[5]), .ZN(n_711));
   AOI22_X1 i_2531 (.A1(in1[22]), .A2(in2[4]), .B1(in1[23]), .B2(in2[3]), 
      .ZN(n_712));
   NAND4_X1 i_2532 (.A1(in1[22]), .A2(in2[4]), .A3(in1[23]), .A4(in2[3]), 
      .ZN(n_713));
   FA_X1 i_2533 (.A(n_3042), .B(n_3035), .CI(n_3028), .CO(n_3089), .S(n_3088));
   FA_X1 i_2534 (.A(n_3063), .B(n_3056), .CI(n_3049), .CO(n_3087), .S(n_3086));
   FA_X1 i_2535 (.A(n_2834), .B(n_2827), .CI(n_2820), .CO(n_2967), .S(n_714));
   FA_X1 i_2536 (.A(n_2967), .B(n_2961), .CI(n_3069), .CO(n_3085), .S(n_715));
   FA_X1 i_2537 (.A(n_3089), .B(n_3087), .CI(n_3085), .CO(n_716), .S(n_3204));
   FA_X1 i_2538 (.A(n_3043), .B(n_3036), .CI(n_3029), .CO(n_717), .S(n_3188));
   FA_X1 i_2539 (.A(n_3064), .B(n_3057), .CI(n_3050), .CO(n_718), .S(n_3186));
   FA_X1 i_2540 (.A(n_3021), .B(n_3014), .CI(n_3005), .CO(n_3091), .S(n_3090));
   FA_X1 i_2541 (.A(n_3188), .B(n_3186), .CI(n_3091), .CO(n_882), .S(n_3202));
   FA_X1 i_2542 (.A(n_3090), .B(n_3088), .CI(n_3086), .CO(n_3101), .S(n_883));
   FA_X1 i_2543 (.A(n_3204), .B(n_3202), .CI(n_3101), .CO(n_885), .S(n_884));
   XNOR2_X1 i_2544 (.A(n_1121), .B(n_886), .ZN(n_3005));
   NOR2_X1 i_2545 (.A1(n_1125), .A2(n_1124), .ZN(n_886));
   XNOR2_X1 i_2546 (.A(n_1178), .B(n_887), .ZN(n_3014));
   NOR2_X1 i_2547 (.A1(n_1181), .A2(n_1180), .ZN(n_887));
   XNOR2_X1 i_2548 (.A(n_1192), .B(n_888), .ZN(n_3021));
   NOR2_X1 i_2549 (.A1(n_1196), .A2(n_1193), .ZN(n_888));
   OAI22_X1 i_2550 (.A1(n_1306), .A2(n_1305), .B1(n_1304), .B2(n_891), .ZN(
      n_3050));
   OAI22_X1 i_2551 (.A1(n_1346), .A2(n_1345), .B1(n_1319), .B2(n_1049), .ZN(
      n_3057));
   OAI22_X1 i_2552 (.A1(n_1351), .A2(n_1350), .B1(n_1347), .B2(n_1080), .ZN(
      n_3064));
   OAI22_X1 i_2553 (.A1(n_1354), .A2(n_1353), .B1(n_1352), .B2(n_1104), .ZN(
      n_3029));
   OAI22_X1 i_2554 (.A1(n_1373), .A2(n_1370), .B1(n_1369), .B2(n_1109), .ZN(
      n_3036));
   OAI22_X1 i_2555 (.A1(n_1376), .A2(n_1375), .B1(n_1374), .B2(n_1112), .ZN(
      n_3043));
   XOR2_X1 i_2556 (.A(n_1199), .B(n_889), .Z(n_3069));
   NAND2_X1 i_2557 (.A1(n_1203), .A2(n_1200), .ZN(n_889));
   AOI21_X1 i_2558 (.A(n_1285), .B1(n_1205), .B2(n_1204), .ZN(n_2961));
   OAI21_X1 i_2559 (.A(n_1291), .B1(n_1290), .B2(n_1289), .ZN(n_2820));
   OAI21_X1 i_2560 (.A(n_1296), .B1(n_1295), .B2(n_1293), .ZN(n_2827));
   OAI21_X1 i_2561 (.A(n_1300), .B1(n_1299), .B2(n_1298), .ZN(n_2834));
   XNOR2_X1 i_2562 (.A(n_1304), .B(n_890), .ZN(n_3049));
   NOR2_X1 i_2563 (.A1(n_892), .A2(n_891), .ZN(n_890));
   AOI22_X1 i_2564 (.A1(in1[22]), .A2(in2[11]), .B1(in1[21]), .B2(in2[12]), 
      .ZN(n_891));
   NOR2_X1 i_2565 (.A1(n_1306), .A2(n_1305), .ZN(n_892));
   XNOR2_X1 i_2566 (.A(n_1319), .B(n_893), .ZN(n_3056));
   NOR2_X1 i_2567 (.A1(n_1050), .A2(n_1049), .ZN(n_893));
   AOI22_X1 i_2568 (.A1(in1[25]), .A2(in2[8]), .B1(in1[24]), .B2(in2[9]), 
      .ZN(n_1049));
   NOR2_X1 i_2569 (.A1(n_1346), .A2(n_1345), .ZN(n_1050));
   XNOR2_X1 i_2570 (.A(n_1347), .B(n_1051), .ZN(n_3063));
   NOR2_X1 i_2571 (.A1(n_1082), .A2(n_1080), .ZN(n_1051));
   AOI22_X1 i_2572 (.A1(in1[28]), .A2(in2[5]), .B1(in1[27]), .B2(in2[6]), 
      .ZN(n_1080));
   NOR2_X1 i_2573 (.A1(n_1351), .A2(n_1350), .ZN(n_1082));
   XNOR2_X1 i_2574 (.A(n_1352), .B(n_1094), .ZN(n_3028));
   NOR2_X1 i_2575 (.A1(n_1105), .A2(n_1104), .ZN(n_1094));
   AOI22_X1 i_2576 (.A1(in1[13]), .A2(in2[20]), .B1(in1[12]), .B2(in2[21]), 
      .ZN(n_1104));
   NOR2_X1 i_2577 (.A1(n_1354), .A2(n_1353), .ZN(n_1105));
   XNOR2_X1 i_2578 (.A(n_1369), .B(n_1106), .ZN(n_3035));
   NOR2_X1 i_2579 (.A1(n_1110), .A2(n_1109), .ZN(n_1106));
   AOI22_X1 i_2580 (.A1(in1[16]), .A2(in2[17]), .B1(in1[15]), .B2(in2[18]), 
      .ZN(n_1109));
   NOR2_X1 i_2581 (.A1(n_1373), .A2(n_1370), .ZN(n_1110));
   XNOR2_X1 i_2582 (.A(n_1374), .B(n_1111), .ZN(n_3042));
   NOR2_X1 i_2583 (.A1(n_1115), .A2(n_1112), .ZN(n_1111));
   AOI22_X1 i_2584 (.A1(in1[19]), .A2(in2[14]), .B1(in1[18]), .B2(in2[15]), 
      .ZN(n_1112));
   NOR2_X1 i_2585 (.A1(n_1376), .A2(n_1375), .ZN(n_1115));
   AND2_X1 i_2586 (.A1(in1[2]), .A2(in2[31]), .ZN(n_1121));
   AOI22_X1 i_2587 (.A1(in1[4]), .A2(in2[29]), .B1(in1[3]), .B2(in2[30]), 
      .ZN(n_1124));
   NOR2_X1 i_2588 (.A1(n_1177), .A2(n_1176), .ZN(n_1125));
   NAND2_X1 i_2589 (.A1(in1[3]), .A2(in2[29]), .ZN(n_1176));
   NAND2_X1 i_2590 (.A1(in1[4]), .A2(in2[30]), .ZN(n_1177));
   NAND2_X1 i_2591 (.A1(in1[5]), .A2(in2[28]), .ZN(n_1178));
   AOI22_X1 i_2592 (.A1(in1[7]), .A2(in2[26]), .B1(in1[6]), .B2(in2[27]), 
      .ZN(n_1180));
   NOR2_X1 i_2593 (.A1(n_1183), .A2(n_1182), .ZN(n_1181));
   NAND2_X1 i_2594 (.A1(in1[6]), .A2(in2[26]), .ZN(n_1182));
   NAND2_X1 i_2595 (.A1(in1[7]), .A2(in2[27]), .ZN(n_1183));
   NAND2_X1 i_2596 (.A1(in1[8]), .A2(in2[25]), .ZN(n_1192));
   AOI22_X1 i_2597 (.A1(in1[10]), .A2(in2[23]), .B1(in1[9]), .B2(in2[24]), 
      .ZN(n_1193));
   NOR2_X1 i_2598 (.A1(n_1198), .A2(n_1197), .ZN(n_1196));
   NAND2_X1 i_2599 (.A1(in1[9]), .A2(in2[23]), .ZN(n_1197));
   NAND2_X1 i_2600 (.A1(in1[10]), .A2(in2[24]), .ZN(n_1198));
   NAND2_X1 i_2601 (.A1(in1[29]), .A2(in2[4]), .ZN(n_1199));
   OAI211_X1 i_2602 (.A(in1[31]), .B(in2[2]), .C1(n_1383), .C2(n_599), .ZN(
      n_1200));
   OAI211_X1 i_2603 (.A(in2[3]), .B(in1[30]), .C1(n_1384), .C2(n_1380), .ZN(
      n_1203));
   OAI211_X1 i_2604 (.A(in1[30]), .B(in2[2]), .C1(n_1384), .C2(n_1377), .ZN(
      n_1204));
   OAI21_X1 i_2605 (.A(n_1206), .B1(n_1212), .B2(n_1210), .ZN(n_1205));
   OAI21_X1 i_2606 (.A(n_1207), .B1(n_1382), .B2(n_1380), .ZN(n_1206));
   NAND2_X1 i_2607 (.A1(in1[28]), .A2(in2[3]), .ZN(n_1207));
   NOR2_X1 i_2608 (.A1(n_1381), .A2(n_693), .ZN(n_1210));
   INV_X1 i_2609 (.A(n_1212), .ZN(n_1211));
   NOR3_X1 i_2610 (.A1(n_1382), .A2(n_1278), .A3(n_599), .ZN(n_1212));
   NAND2_X1 i_2611 (.A1(in1[28]), .A2(in2[2]), .ZN(n_1278));
   INV_X1 i_2612 (.A(n_1286), .ZN(n_1285));
   OAI211_X1 i_2613 (.A(in1[31]), .B(in2[1]), .C1(n_1383), .C2(n_1380), .ZN(
      n_1286));
   NAND2_X1 i_2614 (.A1(in1[18]), .A2(in2[13]), .ZN(n_1289));
   AOI22_X1 i_2615 (.A1(in1[19]), .A2(in2[12]), .B1(in1[20]), .B2(in2[11]), 
      .ZN(n_1290));
   NAND4_X1 i_2616 (.A1(in1[19]), .A2(in2[12]), .A3(in1[20]), .A4(in2[11]), 
      .ZN(n_1291));
   NAND2_X1 i_2617 (.A1(in1[19]), .A2(in2[12]), .ZN(n_1292));
   NAND2_X1 i_2618 (.A1(in1[21]), .A2(in2[10]), .ZN(n_1293));
   AOI22_X1 i_2619 (.A1(in1[22]), .A2(in2[9]), .B1(in1[23]), .B2(in2[8]), 
      .ZN(n_1295));
   NAND4_X1 i_2620 (.A1(in1[22]), .A2(in2[9]), .A3(in1[23]), .A4(in2[8]), 
      .ZN(n_1296));
   NAND2_X1 i_2621 (.A1(in1[22]), .A2(in2[9]), .ZN(n_1297));
   NAND2_X1 i_2622 (.A1(in1[24]), .A2(in2[7]), .ZN(n_1298));
   AOI22_X1 i_2623 (.A1(in1[25]), .A2(in2[6]), .B1(in1[26]), .B2(in2[5]), 
      .ZN(n_1299));
   NAND4_X1 i_2624 (.A1(in1[25]), .A2(in2[6]), .A3(in1[26]), .A4(in2[5]), 
      .ZN(n_1300));
   NAND2_X1 i_2625 (.A1(in1[25]), .A2(in2[6]), .ZN(n_1303));
   NAND2_X1 i_2626 (.A1(in1[20]), .A2(in2[13]), .ZN(n_1304));
   NAND2_X1 i_2627 (.A1(in1[21]), .A2(in2[11]), .ZN(n_1305));
   NAND2_X1 i_2628 (.A1(in1[22]), .A2(in2[12]), .ZN(n_1306));
   NAND2_X1 i_2629 (.A1(in1[23]), .A2(in2[10]), .ZN(n_1319));
   NAND2_X1 i_2630 (.A1(in1[24]), .A2(in2[8]), .ZN(n_1345));
   NAND2_X1 i_2631 (.A1(in1[25]), .A2(in2[9]), .ZN(n_1346));
   NAND2_X1 i_2632 (.A1(in1[26]), .A2(in2[7]), .ZN(n_1347));
   NAND2_X1 i_2633 (.A1(in1[27]), .A2(in2[5]), .ZN(n_1350));
   NAND2_X1 i_2634 (.A1(in1[28]), .A2(in2[6]), .ZN(n_1351));
   NAND2_X1 i_2635 (.A1(in1[11]), .A2(in2[22]), .ZN(n_1352));
   NAND2_X1 i_2636 (.A1(in1[12]), .A2(in2[20]), .ZN(n_1353));
   NAND2_X1 i_2637 (.A1(in1[13]), .A2(in2[21]), .ZN(n_1354));
   NAND2_X1 i_2638 (.A1(in1[14]), .A2(in2[19]), .ZN(n_1369));
   NAND2_X1 i_2639 (.A1(in1[15]), .A2(in2[17]), .ZN(n_1370));
   NAND2_X1 i_2640 (.A1(in1[16]), .A2(in2[18]), .ZN(n_1373));
   NAND2_X1 i_2641 (.A1(in1[17]), .A2(in2[16]), .ZN(n_1374));
   NAND2_X1 i_2642 (.A1(in1[18]), .A2(in2[14]), .ZN(n_1375));
   NAND2_X1 i_2643 (.A1(in1[19]), .A2(in2[15]), .ZN(n_1376));
   INV_X1 i_2644 (.A(in2[1]), .ZN(n_1377));
   INV_X1 i_2645 (.A(in2[2]), .ZN(n_1380));
   INV_X1 i_2646 (.A(in1[27]), .ZN(n_1381));
   INV_X1 i_2647 (.A(in1[29]), .ZN(n_1382));
   INV_X1 i_2648 (.A(in1[30]), .ZN(n_1383));
   INV_X1 i_2649 (.A(in1[31]), .ZN(n_1384));
   FA_X1 i_2650 (.A(n_2792), .B(n_2785), .CI(n_2776), .CO(n_2971), .S(n_2970));
   FA_X1 i_2651 (.A(n_2813), .B(n_2806), .CI(n_2799), .CO(n_2969), .S(n_2968));
   FA_X1 i_2652 (.A(n_1575), .B(n_2971), .CI(n_2969), .CO(n_1387), .S(n_3082));
   FA_X1 i_2653 (.A(n_2805), .B(n_2798), .CI(n_2791), .CO(n_2866), .S(n_1439));
   FA_X1 i_2654 (.A(n_2826), .B(n_2819), .CI(n_2812), .CO(n_2864), .S(n_1440));
   FA_X1 i_2655 (.A(n_714), .B(n_2866), .CI(n_2864), .CO(n_2985), .S(n_1441));
   FA_X1 i_2656 (.A(n_2585), .B(n_2578), .CI(n_2571), .CO(n_2741), .S(n_1442));
   FA_X1 i_2657 (.A(n_2606), .B(n_2599), .CI(n_2592), .CO(n_2739), .S(n_1445));
   FA_X1 i_2658 (.A(n_2741), .B(n_2739), .CI(n_2733), .CO(n_2860), .S(n_1446));
   FA_X1 i_2659 (.A(n_2860), .B(n_2970), .CI(n_2968), .CO(n_2983), .S(n_1447));
   FA_X1 i_2660 (.A(n_3082), .B(n_2985), .CI(n_2983), .CO(n_1449), .S(n_1448));
   AOI21_X1 i_2661 (.A(n_1501), .B1(n_1500), .B2(n_1499), .ZN(n_2733));
   OAI21_X1 i_2662 (.A(n_1519), .B1(n_1518), .B2(n_1517), .ZN(n_2592));
   OAI21_X1 i_2663 (.A(n_1540), .B1(n_1521), .B2(n_1520), .ZN(n_2599));
   OAI21_X1 i_2664 (.A(n_1545), .B1(n_1544), .B2(n_1541), .ZN(n_2606));
   OAI21_X1 i_2665 (.A(n_1548), .B1(n_1547), .B2(n_1546), .ZN(n_2571));
   OAI21_X1 i_2666 (.A(n_1554), .B1(n_1553), .B2(n_1551), .ZN(n_2578));
   OAI21_X1 i_2667 (.A(n_1559), .B1(n_1558), .B2(n_1555), .ZN(n_2585));
   XOR2_X1 i_2668 (.A(n_1487), .B(n_1451), .Z(n_2812));
   OAI21_X1 i_2669 (.A(n_1491), .B1(n_1562), .B2(n_1492), .ZN(n_1451));
   XNOR2_X1 i_2670 (.A(n_1289), .B(n_1452), .ZN(n_2819));
   NOR2_X1 i_2671 (.A1(n_1290), .A2(n_1578), .ZN(n_1452));
   XNOR2_X1 i_2672 (.A(n_1293), .B(n_1455), .ZN(n_2826));
   NOR2_X1 i_2673 (.A1(n_1295), .A2(n_1579), .ZN(n_1455));
   XOR2_X1 i_2674 (.A(n_1493), .B(n_1456), .Z(n_2791));
   OAI21_X1 i_2675 (.A(n_1497), .B1(n_1574), .B2(n_1498), .ZN(n_1456));
   XOR2_X1 i_2676 (.A(n_1461), .B(n_1459), .Z(n_2798));
   OAI21_X1 i_2677 (.A(n_1479), .B1(n_1560), .B2(n_1480), .ZN(n_1459));
   XOR2_X1 i_2678 (.A(n_1483), .B(n_1460), .Z(n_2805));
   OAI21_X1 i_2679 (.A(n_1485), .B1(n_1561), .B2(n_1486), .ZN(n_1460));
   OAI22_X1 i_2680 (.A1(n_1560), .A2(n_1480), .B1(n_1462), .B2(n_1461), .ZN(
      n_2799));
   NAND2_X1 i_2681 (.A1(in2[22]), .A2(in1[9]), .ZN(n_1461));
   INV_X1 i_2682 (.A(n_1479), .ZN(n_1462));
   NAND2_X1 i_2683 (.A1(n_1560), .A2(n_1480), .ZN(n_1479));
   NAND2_X1 i_2684 (.A1(in2[20]), .A2(in1[11]), .ZN(n_1480));
   OAI22_X1 i_2685 (.A1(n_1561), .A2(n_1486), .B1(n_1484), .B2(n_1483), .ZN(
      n_2806));
   NAND2_X1 i_2686 (.A1(in2[19]), .A2(in1[12]), .ZN(n_1483));
   INV_X1 i_2687 (.A(n_1485), .ZN(n_1484));
   NAND2_X1 i_2688 (.A1(n_1561), .A2(n_1486), .ZN(n_1485));
   NAND2_X1 i_2689 (.A1(in2[17]), .A2(in1[14]), .ZN(n_1486));
   OAI22_X1 i_2690 (.A1(n_1562), .A2(n_1492), .B1(n_1490), .B2(n_1487), .ZN(
      n_2813));
   NAND2_X1 i_2691 (.A1(in2[16]), .A2(in1[15]), .ZN(n_1487));
   INV_X1 i_2692 (.A(n_1491), .ZN(n_1490));
   NAND2_X1 i_2693 (.A1(n_1562), .A2(n_1492), .ZN(n_1491));
   NAND2_X1 i_2694 (.A1(in2[14]), .A2(in1[17]), .ZN(n_1492));
   OAI21_X1 i_2695 (.A(n_1567), .B1(n_1566), .B2(n_1565), .ZN(n_2776));
   OAI21_X1 i_2696 (.A(n_1572), .B1(n_1571), .B2(n_1569), .ZN(n_2785));
   OAI22_X1 i_2697 (.A1(n_1574), .A2(n_1498), .B1(n_1494), .B2(n_1493), .ZN(
      n_2792));
   NAND2_X1 i_2698 (.A1(in2[25]), .A2(in1[6]), .ZN(n_1493));
   INV_X1 i_2699 (.A(n_1497), .ZN(n_1494));
   NAND2_X1 i_2700 (.A1(n_1574), .A2(n_1498), .ZN(n_1497));
   NAND2_X1 i_2701 (.A1(in2[23]), .A2(in1[8]), .ZN(n_1498));
   NAND2_X1 i_2702 (.A1(n_1505), .A2(n_1504), .ZN(n_1499));
   NAND2_X1 i_2703 (.A1(in2[0]), .A2(in1[30]), .ZN(n_1500));
   NOR2_X1 i_2704 (.A1(n_1505), .A2(n_1504), .ZN(n_1501));
   OAI21_X1 i_2705 (.A(n_1508), .B1(n_1507), .B2(n_1506), .ZN(n_1504));
   OAI21_X1 i_2706 (.A(n_1513), .B1(n_1512), .B2(n_1511), .ZN(n_1505));
   NAND2_X1 i_2707 (.A1(in2[5]), .A2(in1[24]), .ZN(n_1506));
   AOI22_X1 i_2708 (.A1(in2[3]), .A2(in1[26]), .B1(in2[4]), .B2(in1[25]), 
      .ZN(n_1507));
   NAND4_X1 i_2709 (.A1(in2[3]), .A2(in1[26]), .A3(in2[4]), .A4(in1[25]), 
      .ZN(n_1508));
   NAND2_X1 i_2710 (.A1(in2[2]), .A2(in1[27]), .ZN(n_1511));
   AOI21_X1 i_2711 (.A(n_1514), .B1(in2[0]), .B2(in1[29]), .ZN(n_1512));
   NAND3_X1 i_2712 (.A1(in2[0]), .A2(in1[29]), .A3(n_1514), .ZN(n_1513));
   NOR2_X1 i_2713 (.A1(n_1580), .A2(n_1377), .ZN(n_1514));
   NAND2_X1 i_2714 (.A1(in2[14]), .A2(in1[15]), .ZN(n_1517));
   AOI22_X1 i_2715 (.A1(in2[12]), .A2(in1[17]), .B1(in2[13]), .B2(in1[16]), 
      .ZN(n_1518));
   NAND4_X1 i_2716 (.A1(in2[12]), .A2(in1[17]), .A3(in2[13]), .A4(in1[16]), 
      .ZN(n_1519));
   NAND2_X1 i_2717 (.A1(in2[11]), .A2(in1[18]), .ZN(n_1520));
   AOI22_X1 i_2718 (.A1(in2[9]), .A2(in1[20]), .B1(in2[10]), .B2(in1[19]), 
      .ZN(n_1521));
   NAND4_X1 i_2719 (.A1(in2[9]), .A2(in1[20]), .A3(in2[10]), .A4(in1[19]), 
      .ZN(n_1540));
   NAND2_X1 i_2720 (.A1(in2[8]), .A2(in1[21]), .ZN(n_1541));
   AOI22_X1 i_2721 (.A1(in2[6]), .A2(in1[23]), .B1(in2[7]), .B2(in1[22]), 
      .ZN(n_1544));
   NAND4_X1 i_2722 (.A1(in2[6]), .A2(in1[23]), .A3(in2[7]), .A4(in1[22]), 
      .ZN(n_1545));
   NAND2_X1 i_2723 (.A1(in2[23]), .A2(in1[6]), .ZN(n_1546));
   AOI22_X1 i_2724 (.A1(in2[21]), .A2(in1[8]), .B1(in2[22]), .B2(in1[7]), 
      .ZN(n_1547));
   NAND4_X1 i_2725 (.A1(in2[21]), .A2(in1[8]), .A3(in2[22]), .A4(in1[7]), 
      .ZN(n_1548));
   NAND2_X1 i_2726 (.A1(in2[20]), .A2(in1[9]), .ZN(n_1551));
   AOI22_X1 i_2727 (.A1(in2[18]), .A2(in1[11]), .B1(in2[19]), .B2(in1[10]), 
      .ZN(n_1553));
   NAND4_X1 i_2728 (.A1(in2[18]), .A2(in1[11]), .A3(in2[19]), .A4(in1[10]), 
      .ZN(n_1554));
   NAND2_X1 i_2729 (.A1(in2[17]), .A2(in1[12]), .ZN(n_1555));
   AOI22_X1 i_2730 (.A1(in2[15]), .A2(in1[14]), .B1(in2[16]), .B2(in1[13]), 
      .ZN(n_1558));
   NAND4_X1 i_2731 (.A1(in2[15]), .A2(in1[14]), .A3(in2[16]), .A4(in1[13]), 
      .ZN(n_1559));
   NAND2_X1 i_2732 (.A1(in2[21]), .A2(in1[10]), .ZN(n_1560));
   NAND2_X1 i_2733 (.A1(in2[18]), .A2(in1[13]), .ZN(n_1561));
   NAND2_X1 i_2734 (.A1(in2[15]), .A2(in1[16]), .ZN(n_1562));
   NOR2_X1 i_2735 (.A1(n_1602), .A2(n_690), .ZN(n_1565));
   AOI22_X1 i_2736 (.A1(in2[29]), .A2(in1[2]), .B1(in2[30]), .B2(in1[1]), 
      .ZN(n_1566));
   NAND3_X1 i_2737 (.A1(in2[30]), .A2(in1[2]), .A3(n_1568), .ZN(n_1567));
   NOR2_X1 i_2738 (.A1(n_1581), .A2(n_691), .ZN(n_1568));
   NAND2_X1 i_2739 (.A1(in2[28]), .A2(in1[3]), .ZN(n_1569));
   AOI22_X1 i_2740 (.A1(in2[27]), .A2(in1[4]), .B1(in2[26]), .B2(in1[5]), 
      .ZN(n_1571));
   NAND4_X1 i_2741 (.A1(in2[27]), .A2(in1[4]), .A3(in2[26]), .A4(in1[5]), 
      .ZN(n_1572));
   NAND2_X1 i_2742 (.A1(in2[27]), .A2(in1[4]), .ZN(n_1573));
   NAND2_X1 i_2743 (.A1(in2[24]), .A2(in1[7]), .ZN(n_1574));
   NAND3_X1 i_2744 (.A1(in2[31]), .A2(n_1576), .A3(in1[1]), .ZN(n_1575));
   NAND2_X1 i_2745 (.A1(in2[30]), .A2(in1[2]), .ZN(n_1576));
   INV_X1 i_2746 (.A(n_1291), .ZN(n_1578));
   INV_X1 i_2747 (.A(n_1296), .ZN(n_1579));
   INV_X1 i_2748 (.A(in1[28]), .ZN(n_1580));
   INV_X1 i_2749 (.A(in2[29]), .ZN(n_1581));
   INV_X1 i_2750 (.A(in2[31]), .ZN(n_1602));
   FA_X1 i_2751 (.A(n_3138), .B(n_3131), .CI(n_3124), .CO(n_3199), .S(n_3198));
   FA_X1 i_2752 (.A(n_3159), .B(n_3152), .CI(n_3145), .CO(n_3197), .S(n_3196));
   FA_X1 i_2753 (.A(n_3180), .B(n_3173), .CI(n_3166), .CO(n_3195), .S(n_3194));
   FA_X1 i_2754 (.A(n_3199), .B(n_3197), .CI(n_3195), .CO(n_1603), .S(n_3304));
   FA_X1 i_2755 (.A(n_3139), .B(n_3132), .CI(n_3125), .CO(n_1606), .S(n_3290));
   FA_X1 i_2756 (.A(n_3160), .B(n_3153), .CI(n_3146), .CO(n_1607), .S(n_3288));
   FA_X1 i_2757 (.A(n_541), .B(n_3174), .CI(n_3167), .CO(n_1608), .S(n_3286));
   FA_X1 i_2758 (.A(n_3290), .B(n_3288), .CI(n_3286), .CO(n_1609), .S(n_3302));
   FA_X1 i_2759 (.A(n_3198), .B(n_3196), .CI(n_3194), .CO(n_3209), .S(n_1610));
   FA_X1 i_2760 (.A(n_3304), .B(n_3302), .CI(n_3209), .CO(n_1614), .S(n_1613));
   OAI22_X1 i_2761 (.A1(n_1346), .A2(n_1620), .B1(n_1617), .B2(n_1615), .ZN(
      n_3167));
   OAI22_X1 i_2762 (.A1(n_1351), .A2(n_1624), .B1(n_1623), .B2(n_1621), .ZN(
      n_3174));
   NAND2_X1 i_2763 (.A1(in2[4]), .A2(in1[31]), .ZN(n_541));
   OAI22_X1 i_2764 (.A1(n_1373), .A2(n_1630), .B1(n_1629), .B2(n_1627), .ZN(
      n_3146));
   OAI22_X1 i_2765 (.A1(n_1376), .A2(n_1636), .B1(n_1635), .B2(n_1631), .ZN(
      n_3153));
   OAI22_X1 i_2766 (.A1(n_1306), .A2(n_1641), .B1(n_1640), .B2(n_1637), .ZN(
      n_3160));
   OAI22_X1 i_2767 (.A1(n_1183), .A2(n_1645), .B1(n_1644), .B2(n_1642), .ZN(
      n_3125));
   OAI22_X1 i_2768 (.A1(n_1198), .A2(n_1651), .B1(n_1650), .B2(n_1648), .ZN(
      n_3132));
   OAI22_X1 i_2769 (.A1(n_1354), .A2(n_1677), .B1(n_1676), .B2(n_1672), .ZN(
      n_3139));
   XNOR2_X1 i_2770 (.A(n_1616), .B(n_1615), .ZN(n_3166));
   NAND2_X1 i_2771 (.A1(in2[10]), .A2(in1[24]), .ZN(n_1615));
   XOR2_X1 i_2772 (.A(n_1346), .B(n_1620), .Z(n_1616));
   AND2_X1 i_2773 (.A1(n_1346), .A2(n_1620), .ZN(n_1617));
   NAND2_X1 i_2774 (.A1(in2[8]), .A2(in1[26]), .ZN(n_1620));
   XNOR2_X1 i_2775 (.A(n_1622), .B(n_1621), .ZN(n_3173));
   NAND2_X1 i_2776 (.A1(in2[7]), .A2(in1[27]), .ZN(n_1621));
   XOR2_X1 i_2777 (.A(n_1351), .B(n_1624), .Z(n_1622));
   AND2_X1 i_2778 (.A1(n_1351), .A2(n_1624), .ZN(n_1623));
   NAND2_X1 i_2779 (.A1(in2[5]), .A2(in1[29]), .ZN(n_1624));
   XNOR2_X1 i_2780 (.A(n_1679), .B(n_1678), .ZN(n_3180));
   XNOR2_X1 i_2781 (.A(n_1628), .B(n_1627), .ZN(n_3145));
   NAND2_X1 i_2782 (.A1(in2[19]), .A2(in1[15]), .ZN(n_1627));
   XOR2_X1 i_2783 (.A(n_1373), .B(n_1630), .Z(n_1628));
   AND2_X1 i_2784 (.A1(n_1373), .A2(n_1630), .ZN(n_1629));
   NAND2_X1 i_2785 (.A1(in2[17]), .A2(in1[17]), .ZN(n_1630));
   XNOR2_X1 i_2786 (.A(n_1634), .B(n_1631), .ZN(n_3152));
   NAND2_X1 i_2787 (.A1(in2[16]), .A2(in1[18]), .ZN(n_1631));
   XOR2_X1 i_2788 (.A(n_1376), .B(n_1636), .Z(n_1634));
   AND2_X1 i_2789 (.A1(n_1376), .A2(n_1636), .ZN(n_1635));
   NAND2_X1 i_2790 (.A1(in2[14]), .A2(in1[20]), .ZN(n_1636));
   XNOR2_X1 i_2791 (.A(n_1638), .B(n_1637), .ZN(n_3159));
   NAND2_X1 i_2792 (.A1(in2[13]), .A2(in1[21]), .ZN(n_1637));
   XOR2_X1 i_2793 (.A(n_1306), .B(n_1641), .Z(n_1638));
   AND2_X1 i_2794 (.A1(n_1306), .A2(n_1641), .ZN(n_1640));
   NAND2_X1 i_2795 (.A1(in2[11]), .A2(in1[23]), .ZN(n_1641));
   XNOR2_X1 i_2796 (.A(n_1643), .B(n_1642), .ZN(n_3124));
   NAND2_X1 i_2797 (.A1(in2[28]), .A2(in1[6]), .ZN(n_1642));
   XOR2_X1 i_2798 (.A(n_1183), .B(n_1645), .Z(n_1643));
   AND2_X1 i_2799 (.A1(n_1183), .A2(n_1645), .ZN(n_1644));
   NAND2_X1 i_2800 (.A1(in2[26]), .A2(in1[8]), .ZN(n_1645));
   XNOR2_X1 i_2801 (.A(n_1649), .B(n_1648), .ZN(n_3131));
   NAND2_X1 i_2802 (.A1(in2[25]), .A2(in1[9]), .ZN(n_1648));
   XOR2_X1 i_2803 (.A(n_1198), .B(n_1651), .Z(n_1649));
   AND2_X1 i_2804 (.A1(n_1198), .A2(n_1651), .ZN(n_1650));
   NAND2_X1 i_2805 (.A1(in2[23]), .A2(in1[11]), .ZN(n_1651));
   XNOR2_X1 i_2806 (.A(n_1673), .B(n_1672), .ZN(n_3138));
   NAND2_X1 i_2807 (.A1(in2[22]), .A2(in1[12]), .ZN(n_1672));
   XOR2_X1 i_2808 (.A(n_1354), .B(n_1677), .Z(n_1673));
   AND2_X1 i_2809 (.A1(n_1354), .A2(n_1677), .ZN(n_1676));
   NAND2_X1 i_2810 (.A1(in2[20]), .A2(in1[14]), .ZN(n_1677));
   OAI21_X1 i_2811 (.A(n_1203), .B1(n_1684), .B2(n_1199), .ZN(n_1678));
   XOR2_X1 i_2812 (.A(n_1683), .B(n_1680), .Z(n_1679));
   NOR2_X1 i_2813 (.A1(n_1384), .A2(n_599), .ZN(n_1680));
   NOR2_X1 i_2814 (.A1(n_1383), .A2(n_693), .ZN(n_1683));
   INV_X1 i_2815 (.A(n_1200), .ZN(n_1684));
   FA_X1 i_2816 (.A(n_2912), .B(n_2905), .CI(n_2898), .CO(n_3081), .S(n_3080));
   FA_X1 i_2817 (.A(n_2933), .B(n_2926), .CI(n_2919), .CO(n_3079), .S(n_3078));
   FA_X1 i_2818 (.A(n_2954), .B(n_2947), .CI(n_2940), .CO(n_3077), .S(n_3076));
   FA_X1 i_2819 (.A(n_3081), .B(n_3079), .CI(n_3077), .CO(n_1685), .S(n_3192));
   FA_X1 i_2820 (.A(n_2904), .B(n_2897), .CI(n_2892), .CO(n_2981), .S(n_1686));
   FA_X1 i_2821 (.A(n_2925), .B(n_2918), .CI(n_2911), .CO(n_2979), .S(n_1687));
   FA_X1 i_2822 (.A(n_3076), .B(n_2981), .CI(n_2979), .CO(n_3095), .S(n_1690));
   FA_X1 i_2823 (.A(n_2677), .B(n_2670), .CI(n_2663), .CO(n_2858), .S(n_1691));
   FA_X1 i_2824 (.A(n_2698), .B(n_2691), .CI(n_2684), .CO(n_2856), .S(n_1692));
   FA_X1 i_2825 (.A(n_2719), .B(n_2712), .CI(n_2705), .CO(n_2854), .S(n_1693));
   FA_X1 i_2826 (.A(n_2858), .B(n_2856), .CI(n_2854), .CO(n_2973), .S(n_1694));
   FA_X1 i_2827 (.A(n_2973), .B(n_3080), .CI(n_3078), .CO(n_3093), .S(n_1697));
   FA_X1 i_2828 (.A(n_3192), .B(n_3095), .CI(n_3093), .CO(n_1699), .S(n_1698));
   OAI21_X1 i_2829 (.A(n_1748), .B1(n_1745), .B2(n_1744), .ZN(n_2705));
   OAI21_X1 i_2830 (.A(n_1751), .B1(n_1750), .B2(n_1749), .ZN(n_2712));
   OAI21_X1 i_2831 (.A(n_1756), .B1(n_1755), .B2(n_1752), .ZN(n_2719));
   OAI21_X1 i_2832 (.A(n_1759), .B1(n_1758), .B2(n_1757), .ZN(n_2684));
   OAI21_X1 i_2833 (.A(n_1764), .B1(n_1763), .B2(n_1762), .ZN(n_2691));
   OAI21_X1 i_2834 (.A(n_1769), .B1(n_1766), .B2(n_1765), .ZN(n_2698));
   OAI21_X1 i_2835 (.A(n_1772), .B1(n_1771), .B2(n_1770), .ZN(n_2663));
   OAI21_X1 i_2836 (.A(n_1777), .B1(n_1776), .B2(n_1773), .ZN(n_2670));
   OAI21_X1 i_2837 (.A(n_1780), .B1(n_1779), .B2(n_1778), .ZN(n_2677));
   XOR2_X1 i_2838 (.A(n_1197), .B(n_1700), .Z(n_2911));
   OAI21_X1 i_2839 (.A(n_1720), .B1(n_1352), .B2(n_1560), .ZN(n_1700));
   XOR2_X1 i_2840 (.A(n_1353), .B(n_1701), .Z(n_2918));
   OAI21_X1 i_2841 (.A(n_1708), .B1(n_1369), .B2(n_1561), .ZN(n_1701));
   XOR2_X1 i_2842 (.A(n_1370), .B(n_1704), .Z(n_2925));
   OAI21_X1 i_2843 (.A(n_1712), .B1(n_1374), .B2(n_1562), .ZN(n_1704));
   OAI21_X1 i_2844 (.A(n_1575), .B1(n_1576), .B2(n_1705), .ZN(n_2892));
   NOR2_X1 i_2845 (.A1(n_1602), .A2(n_691), .ZN(n_1705));
   XOR2_X1 i_2846 (.A(n_1176), .B(n_1706), .Z(n_2897));
   OAI21_X1 i_2847 (.A(n_1714), .B1(n_1178), .B2(n_1573), .ZN(n_1706));
   XOR2_X1 i_2848 (.A(n_1182), .B(n_1707), .Z(n_2904));
   OAI21_X1 i_2849 (.A(n_1718), .B1(n_1192), .B2(n_1574), .ZN(n_1707));
   OAI22_X1 i_2850 (.A1(n_1319), .A2(n_1297), .B1(n_1305), .B2(n_1782), .ZN(
      n_2940));
   OAI22_X1 i_2851 (.A1(n_1347), .A2(n_1303), .B1(n_1345), .B2(n_1824), .ZN(
      n_2947));
   OAI22_X1 i_2852 (.A1(n_1199), .A2(n_1207), .B1(n_1350), .B2(n_1828), .ZN(
      n_2954));
   OAI22_X1 i_2853 (.A1(n_1369), .A2(n_1561), .B1(n_1353), .B2(n_1711), .ZN(
      n_2919));
   INV_X1 i_2854 (.A(n_1711), .ZN(n_1708));
   AOI22_X1 i_2855 (.A1(in2[18]), .A2(in1[14]), .B1(in2[19]), .B2(in1[13]), 
      .ZN(n_1711));
   OAI22_X1 i_2856 (.A1(n_1374), .A2(n_1562), .B1(n_1370), .B2(n_1713), .ZN(
      n_2926));
   INV_X1 i_2857 (.A(n_1713), .ZN(n_1712));
   AOI22_X1 i_2858 (.A1(in2[15]), .A2(in1[17]), .B1(in2[16]), .B2(in1[16]), 
      .ZN(n_1713));
   OAI22_X1 i_2859 (.A1(n_1304), .A2(n_1292), .B1(n_1375), .B2(n_1830), .ZN(
      n_2933));
   OAI22_X1 i_2860 (.A1(n_1178), .A2(n_1573), .B1(n_1176), .B2(n_1717), .ZN(
      n_2898));
   INV_X1 i_2861 (.A(n_1717), .ZN(n_1714));
   AOI22_X1 i_2862 (.A1(in2[27]), .A2(in1[5]), .B1(in2[28]), .B2(in1[4]), 
      .ZN(n_1717));
   OAI22_X1 i_2863 (.A1(n_1192), .A2(n_1574), .B1(n_1182), .B2(n_1719), .ZN(
      n_2905));
   INV_X1 i_2864 (.A(n_1719), .ZN(n_1718));
   AOI22_X1 i_2865 (.A1(in2[24]), .A2(in1[8]), .B1(in2[25]), .B2(in1[7]), 
      .ZN(n_1719));
   OAI22_X1 i_2866 (.A1(n_1352), .A2(n_1560), .B1(n_1197), .B2(n_1721), .ZN(
      n_2912));
   INV_X1 i_2867 (.A(n_1721), .ZN(n_1720));
   AOI22_X1 i_2868 (.A1(in2[21]), .A2(in1[11]), .B1(in2[22]), .B2(in1[10]), 
      .ZN(n_1721));
   NAND2_X1 i_2869 (.A1(in2[12]), .A2(in1[18]), .ZN(n_1744));
   AOI22_X1 i_2870 (.A1(in2[10]), .A2(in1[20]), .B1(in2[11]), .B2(in1[19]), 
      .ZN(n_1745));
   NAND4_X1 i_2871 (.A1(in2[10]), .A2(in1[20]), .A3(in2[11]), .A4(in1[19]), 
      .ZN(n_1748));
   NAND2_X1 i_2872 (.A1(in2[9]), .A2(in1[21]), .ZN(n_1749));
   AOI22_X1 i_2873 (.A1(in2[7]), .A2(in1[23]), .B1(in2[8]), .B2(in1[22]), 
      .ZN(n_1750));
   NAND4_X1 i_2874 (.A1(in2[7]), .A2(in1[23]), .A3(in2[8]), .A4(in1[22]), 
      .ZN(n_1751));
   NAND2_X1 i_2875 (.A1(in2[6]), .A2(in1[24]), .ZN(n_1752));
   AOI22_X1 i_2876 (.A1(in2[4]), .A2(in1[26]), .B1(in2[5]), .B2(in1[25]), 
      .ZN(n_1755));
   NAND4_X1 i_2877 (.A1(in2[4]), .A2(in1[26]), .A3(in2[5]), .A4(in1[25]), 
      .ZN(n_1756));
   NAND2_X1 i_2878 (.A1(in2[21]), .A2(in1[9]), .ZN(n_1757));
   AOI22_X1 i_2879 (.A1(in2[19]), .A2(in1[11]), .B1(in2[20]), .B2(in1[10]), 
      .ZN(n_1758));
   NAND4_X1 i_2880 (.A1(in2[19]), .A2(in1[11]), .A3(in2[20]), .A4(in1[10]), 
      .ZN(n_1759));
   NAND2_X1 i_2881 (.A1(in2[18]), .A2(in1[12]), .ZN(n_1762));
   AOI22_X1 i_2882 (.A1(in2[16]), .A2(in1[14]), .B1(in2[17]), .B2(in1[13]), 
      .ZN(n_1763));
   NAND4_X1 i_2883 (.A1(in2[16]), .A2(in1[14]), .A3(in2[17]), .A4(in1[13]), 
      .ZN(n_1764));
   NAND2_X1 i_2884 (.A1(in2[15]), .A2(in1[15]), .ZN(n_1765));
   AOI22_X1 i_2885 (.A1(in2[13]), .A2(in1[17]), .B1(in2[14]), .B2(in1[16]), 
      .ZN(n_1766));
   NAND4_X1 i_2886 (.A1(in2[13]), .A2(in1[17]), .A3(in2[14]), .A4(in1[16]), 
      .ZN(n_1769));
   NAND2_X1 i_2887 (.A1(in2[30]), .A2(in1[0]), .ZN(n_1770));
   AOI21_X1 i_2888 (.A(n_1568), .B1(in2[28]), .B2(in1[2]), .ZN(n_1771));
   NAND3_X1 i_2889 (.A1(in2[28]), .A2(n_1568), .A3(in1[2]), .ZN(n_1772));
   NAND2_X1 i_2890 (.A1(in2[27]), .A2(in1[3]), .ZN(n_1773));
   AOI22_X1 i_2891 (.A1(in2[25]), .A2(in1[5]), .B1(in2[26]), .B2(in1[4]), 
      .ZN(n_1776));
   NAND4_X1 i_2892 (.A1(in2[25]), .A2(in1[5]), .A3(in2[26]), .A4(in1[4]), 
      .ZN(n_1777));
   NAND2_X1 i_2893 (.A1(in2[24]), .A2(in1[6]), .ZN(n_1778));
   AOI22_X1 i_2894 (.A1(in2[22]), .A2(in1[8]), .B1(in2[23]), .B2(in1[7]), 
      .ZN(n_1779));
   NAND4_X1 i_2895 (.A1(in2[22]), .A2(in1[8]), .A3(in2[23]), .A4(in1[7]), 
      .ZN(n_1780));
   AOI22_X1 i_2896 (.A1(in2[9]), .A2(in1[23]), .B1(in2[10]), .B2(in1[22]), 
      .ZN(n_1782));
   NOR2_X1 i_2897 (.A1(n_1319), .A2(n_1297), .ZN(n_1791));
   AOI22_X1 i_2898 (.A1(in2[6]), .A2(in1[26]), .B1(in2[7]), .B2(in1[25]), 
      .ZN(n_1824));
   NOR2_X1 i_2899 (.A1(n_1347), .A2(n_1303), .ZN(n_1825));
   AOI22_X1 i_2900 (.A1(in2[4]), .A2(in1[28]), .B1(in2[3]), .B2(in1[29]), 
      .ZN(n_1828));
   NOR2_X1 i_2901 (.A1(n_1199), .A2(n_1207), .ZN(n_1829));
   AOI22_X1 i_2902 (.A1(in2[12]), .A2(in1[20]), .B1(in2[13]), .B2(in1[19]), 
      .ZN(n_1830));
   NOR2_X1 i_2903 (.A1(n_1304), .A2(n_1292), .ZN(n_1831));
   FA_X1 i_2904 (.A(n_3022), .B(n_3015), .CI(n_3006), .CO(n_3191), .S(n_1832));
   FA_X1 i_2905 (.A(n_3116), .B(n_3191), .CI(n_717), .CO(n_3293), .S(n_1835));
   FA_X1 i_2906 (.A(n_3240), .B(n_3233), .CI(n_3224), .CO(n_1836), .S(n_3391));
   FA_X1 i_2907 (.A(n_3261), .B(n_3254), .CI(n_3247), .CO(n_1837), .S(n_3389));
   FA_X1 i_2908 (.A(n_3293), .B(n_3391), .CI(n_3389), .CO(n_1839), .S(n_1838));
   NAND4_X1 i_2909 (.A1(in2[21]), .A2(in1[14]), .A3(in2[20]), .A4(in1[15]), 
      .ZN(n_1842));
   AOI22_X1 i_2910 (.A1(in2[21]), .A2(in1[14]), .B1(in2[20]), .B2(in1[15]), 
      .ZN(n_1843));
   NAND2_X1 i_2911 (.A1(in2[22]), .A2(in1[13]), .ZN(n_1844));
   OAI21_X1 i_2912 (.A(n_1842), .B1(n_1843), .B2(n_1844), .ZN(n_3247));
   NAND4_X1 i_2913 (.A1(in2[18]), .A2(in1[17]), .A3(in2[17]), .A4(in1[18]), 
      .ZN(n_1845));
   AOI22_X1 i_2914 (.A1(in2[18]), .A2(in1[17]), .B1(in2[17]), .B2(in1[18]), 
      .ZN(n_1846));
   NAND2_X1 i_2915 (.A1(in2[19]), .A2(in1[16]), .ZN(n_1849));
   OAI21_X1 i_2916 (.A(n_1845), .B1(n_1846), .B2(n_1849), .ZN(n_3254));
   NAND4_X1 i_2917 (.A1(in2[15]), .A2(in1[20]), .A3(in2[14]), .A4(in1[21]), 
      .ZN(n_1850));
   AOI22_X1 i_2918 (.A1(in2[15]), .A2(in1[20]), .B1(in2[14]), .B2(in1[21]), 
      .ZN(n_1851));
   NAND2_X1 i_2919 (.A1(in2[16]), .A2(in1[19]), .ZN(n_1852));
   OAI21_X1 i_2920 (.A(n_1850), .B1(n_1851), .B2(n_1852), .ZN(n_3261));
   NAND4_X1 i_2921 (.A1(in2[30]), .A2(in1[6]), .A3(in2[29]), .A4(in1[5]), 
      .ZN(n_1853));
   AOI22_X1 i_2922 (.A1(in2[30]), .A2(in1[5]), .B1(in1[6]), .B2(in2[29]), 
      .ZN(n_1856));
   INV_X1 i_2923 (.A(in1[4]), .ZN(n_1857));
   NOR2_X1 i_2924 (.A1(n_1857), .A2(n_1602), .ZN(n_1858));
   OAI21_X1 i_2925 (.A(n_1853), .B1(n_1856), .B2(n_1858), .ZN(n_3224));
   NAND4_X1 i_2926 (.A1(in2[27]), .A2(in1[8]), .A3(in2[26]), .A4(in1[9]), 
      .ZN(n_1859));
   AOI22_X1 i_2927 (.A1(in2[27]), .A2(in1[8]), .B1(in2[26]), .B2(in1[9]), 
      .ZN(n_1860));
   NAND2_X1 i_2928 (.A1(in2[28]), .A2(in1[7]), .ZN(n_1862));
   OAI21_X1 i_2929 (.A(n_1859), .B1(n_1860), .B2(n_1862), .ZN(n_3233));
   NAND4_X1 i_2930 (.A1(in2[24]), .A2(in1[11]), .A3(in2[23]), .A4(in1[12]), 
      .ZN(n_1863));
   AOI22_X1 i_2931 (.A1(in2[24]), .A2(in1[11]), .B1(in2[23]), .B2(in1[12]), 
      .ZN(n_1864));
   NAND2_X1 i_2932 (.A1(in2[25]), .A2(in1[10]), .ZN(n_1865));
   OAI21_X1 i_2933 (.A(n_1863), .B1(n_1864), .B2(n_1865), .ZN(n_3240));
   INV_X1 i_2934 (.A(n_1125), .ZN(n_1866));
   AOI21_X1 i_2935 (.A(n_1124), .B1(n_1866), .B2(n_1121), .ZN(n_3006));
   INV_X1 i_2936 (.A(n_1181), .ZN(n_1867));
   OAI21_X1 i_2937 (.A(n_1867), .B1(n_1180), .B2(n_1178), .ZN(n_3015));
   INV_X1 i_2938 (.A(n_1196), .ZN(n_1870));
   OAI21_X1 i_2939 (.A(n_1870), .B1(n_1193), .B2(n_1192), .ZN(n_3022));
   INV_X1 i_2940 (.A(n_1177), .ZN(n_1871));
   NAND3_X1 i_2941 (.A1(n_1871), .A2(in2[29]), .A3(in1[5]), .ZN(n_1872));
   AOI21_X1 i_2942 (.A(n_1871), .B1(in2[29]), .B2(in1[5]), .ZN(n_1903));
   INV_X1 i_2943 (.A(n_1903), .ZN(n_1904));
   AND2_X1 i_2944 (.A1(in2[31]), .A2(in1[3]), .ZN(n_1905));
   OAI21_X1 i_2945 (.A(n_1872), .B1(n_1905), .B2(n_1903), .ZN(n_3116));
   FA_X1 i_2946 (.A(n_3354), .B(n_3347), .CI(n_3340), .CO(n_3489), .S(n_1906));
   FA_X1 i_2947 (.A(n_3375), .B(n_3368), .CI(n_3361), .CO(n_3487), .S(n_1909));
   FA_X1 i_2948 (.A(n_3489), .B(n_3487), .CI(n_3481), .CO(n_3582), .S(n_1910));
   FA_X1 i_2949 (.A(n_3439), .B(n_3432), .CI(n_3423), .CO(n_3580), .S(n_1911));
   FA_X1 i_2950 (.A(n_3529), .B(n_3520), .CI(n_3580), .CO(n_1912), .S(n_3669));
   FA_X1 i_2951 (.A(n_3608), .B(n_3582), .CI(n_3669), .CO(n_1916), .S(n_1913));
   OAI21_X1 i_2952 (.A(n_1927), .B1(n_1926), .B2(n_1925), .ZN(n_3423));
   OAI21_X1 i_2953 (.A(n_1932), .B1(n_1931), .B2(n_1930), .ZN(n_3432));
   OAI21_X1 i_2954 (.A(n_1937), .B1(n_1934), .B2(n_1933), .ZN(n_3439));
   AOI21_X1 i_2955 (.A(n_1940), .B1(n_1941), .B2(n_1939), .ZN(n_3520));
   OAI21_X1 i_2956 (.A(n_1946), .B1(n_1945), .B2(n_1944), .ZN(n_3529));
   OAI21_X1 i_2957 (.A(n_1917), .B1(n_1952), .B2(n_1951), .ZN(n_3481));
   NAND2_X1 i_2958 (.A1(n_1953), .A2(n_1950), .ZN(n_1917));
   OAI21_X1 i_2959 (.A(n_1988), .B1(n_1987), .B2(n_1986), .ZN(n_3361));
   OAI21_X1 i_2960 (.A(n_1993), .B1(n_1992), .B2(n_1989), .ZN(n_3368));
   OAI21_X1 i_2961 (.A(n_1996), .B1(n_1995), .B2(n_1994), .ZN(n_3375));
   OAI21_X1 i_2962 (.A(n_2001), .B1(n_2000), .B2(n_1999), .ZN(n_3340));
   OAI21_X1 i_2963 (.A(n_2070), .B1(n_2003), .B2(n_2002), .ZN(n_3347));
   OAI21_X1 i_2964 (.A(n_2073), .B1(n_2072), .B2(n_2071), .ZN(n_3354));
   XNOR2_X1 i_2965 (.A(n_2076), .B(n_1918), .ZN(n_3608));
   AOI21_X1 i_2966 (.A(n_2078), .B1(n_2080), .B2(n_2079), .ZN(n_1918));
   AND2_X1 i_2967 (.A1(in2[31]), .A2(in1[6]), .ZN(n_1925));
   AOI22_X1 i_2968 (.A1(in2[29]), .A2(in1[8]), .B1(in2[30]), .B2(in1[7]), 
      .ZN(n_1926));
   NAND4_X1 i_2969 (.A1(in2[30]), .A2(in2[29]), .A3(in1[8]), .A4(in1[7]), 
      .ZN(n_1927));
   NAND2_X1 i_2970 (.A1(in2[28]), .A2(in1[9]), .ZN(n_1930));
   AOI22_X1 i_2971 (.A1(in2[26]), .A2(in1[11]), .B1(in2[27]), .B2(in1[10]), 
      .ZN(n_1931));
   NAND4_X1 i_2972 (.A1(in2[26]), .A2(in1[11]), .A3(in2[27]), .A4(in1[10]), 
      .ZN(n_1932));
   NAND2_X1 i_2973 (.A1(in2[25]), .A2(in1[12]), .ZN(n_1933));
   AOI21_X1 i_2974 (.A(n_1938), .B1(in2[24]), .B2(in1[13]), .ZN(n_1934));
   NAND3_X1 i_2975 (.A1(in2[24]), .A2(in1[13]), .A3(n_1938), .ZN(n_1937));
   AND2_X1 i_2976 (.A1(in2[23]), .A2(in1[14]), .ZN(n_1938));
   AND2_X1 i_2977 (.A1(in2[31]), .A2(in1[7]), .ZN(n_1939));
   AOI22_X1 i_2978 (.A1(in2[30]), .A2(in1[8]), .B1(in2[29]), .B2(in1[9]), 
      .ZN(n_1940));
   NAND3_X1 i_2979 (.A1(in2[29]), .A2(in1[8]), .A3(n_2080), .ZN(n_1941));
   NAND2_X1 i_2980 (.A1(in2[28]), .A2(in1[10]), .ZN(n_1944));
   AOI22_X1 i_2981 (.A1(in2[27]), .A2(in1[11]), .B1(in2[26]), .B2(in1[12]), 
      .ZN(n_1945));
   NAND4_X1 i_2982 (.A1(in2[26]), .A2(in1[11]), .A3(in2[27]), .A4(in1[12]), 
      .ZN(n_1946));
   OAI21_X1 i_2983 (.A(n_1950), .B1(n_1952), .B2(n_1951), .ZN(n_1947));
   NAND2_X1 i_2984 (.A1(n_1952), .A2(n_1951), .ZN(n_1950));
   NOR2_X1 i_2985 (.A1(n_2083), .A2(n_1384), .ZN(n_1951));
   NAND2_X1 i_2986 (.A1(in2[7]), .A2(in1[30]), .ZN(n_1952));
   OAI21_X1 i_2987 (.A(n_1985), .B1(n_1981), .B2(n_1954), .ZN(n_1953));
   NAND2_X1 i_2988 (.A1(in2[7]), .A2(in1[29]), .ZN(n_1954));
   INV_X1 i_2989 (.A(n_1982), .ZN(n_1981));
   OAI211_X1 i_2990 (.A(in2[5]), .B(in1[31]), .C1(n_2083), .C2(n_1383), .ZN(
      n_1982));
   OAI211_X1 i_2991 (.A(in2[6]), .B(in1[30]), .C1(n_1384), .C2(n_694), .ZN(
      n_1985));
   NAND2_X1 i_2992 (.A1(in2[16]), .A2(in1[20]), .ZN(n_1986));
   AOI22_X1 i_2993 (.A1(in2[15]), .A2(in1[21]), .B1(in2[14]), .B2(in1[22]), 
      .ZN(n_1987));
   NAND4_X1 i_2994 (.A1(in2[15]), .A2(in1[21]), .A3(in2[14]), .A4(in1[22]), 
      .ZN(n_1988));
   NAND2_X1 i_2995 (.A1(in2[13]), .A2(in1[23]), .ZN(n_1989));
   AOI22_X1 i_2996 (.A1(in2[12]), .A2(in1[24]), .B1(in2[11]), .B2(in1[25]), 
      .ZN(n_1992));
   NAND4_X1 i_2997 (.A1(in2[12]), .A2(in1[24]), .A3(in2[11]), .A4(in1[25]), 
      .ZN(n_1993));
   NAND2_X1 i_2998 (.A1(in2[10]), .A2(in1[26]), .ZN(n_1994));
   AOI22_X1 i_2999 (.A1(in2[9]), .A2(in1[27]), .B1(in2[8]), .B2(in1[28]), 
      .ZN(n_1995));
   NAND4_X1 i_3000 (.A1(in2[9]), .A2(in1[27]), .A3(in2[8]), .A4(in1[28]), 
      .ZN(n_1996));
   NAND2_X1 i_3001 (.A1(in2[25]), .A2(in1[11]), .ZN(n_1999));
   AOI22_X1 i_3002 (.A1(in2[24]), .A2(in1[12]), .B1(in2[23]), .B2(in1[13]), 
      .ZN(n_2000));
   NAND4_X1 i_3003 (.A1(in2[24]), .A2(in1[12]), .A3(in2[23]), .A4(in1[13]), 
      .ZN(n_2001));
   NAND2_X1 i_3004 (.A1(in2[22]), .A2(in1[14]), .ZN(n_2002));
   AOI22_X1 i_3005 (.A1(in2[21]), .A2(in1[15]), .B1(in2[20]), .B2(in1[16]), 
      .ZN(n_2003));
   NAND4_X1 i_3006 (.A1(in2[21]), .A2(in1[15]), .A3(in2[20]), .A4(in1[16]), 
      .ZN(n_2070));
   NAND2_X1 i_3007 (.A1(in2[19]), .A2(in1[17]), .ZN(n_2071));
   AOI22_X1 i_3008 (.A1(in2[18]), .A2(in1[18]), .B1(in2[17]), .B2(in1[19]), 
      .ZN(n_2072));
   NAND4_X1 i_3009 (.A1(in2[18]), .A2(in1[18]), .A3(in2[17]), .A4(in1[19]), 
      .ZN(n_2073));
   AND2_X1 i_3010 (.A1(in2[31]), .A2(in1[8]), .ZN(n_2076));
   NAND2_X1 i_3011 (.A1(n_2080), .A2(n_2079), .ZN(n_2077));
   NOR2_X1 i_3012 (.A1(n_2080), .A2(n_2079), .ZN(n_2078));
   AND2_X1 i_3013 (.A1(in2[29]), .A2(in1[10]), .ZN(n_2079));
   AND2_X1 i_3014 (.A1(in2[30]), .A2(in1[9]), .ZN(n_2080));
   INV_X1 i_3015 (.A(in2[6]), .ZN(n_2083));
   OAI21_X1 i_3016 (.A(n_2085), .B1(n_2091), .B2(n_2090), .ZN(n_2084));
   NAND2_X1 i_3017 (.A1(n_2092), .A2(n_2087), .ZN(n_2085));
   OAI21_X1 i_3018 (.A(n_2087), .B1(n_2091), .B2(n_2090), .ZN(n_2086));
   NAND2_X1 i_3019 (.A1(n_2091), .A2(n_2090), .ZN(n_2087));
   NOR2_X1 i_3020 (.A1(n_2262), .A2(n_1384), .ZN(n_2090));
   NAND2_X1 i_3021 (.A1(in1[30]), .A2(in2[13]), .ZN(n_2091));
   OAI21_X1 i_3022 (.A(n_2258), .B1(n_2256), .B2(n_2093), .ZN(n_2092));
   NAND2_X1 i_3023 (.A1(in1[29]), .A2(in2[13]), .ZN(n_2093));
   INV_X1 i_3024 (.A(n_2257), .ZN(n_2256));
   OAI211_X1 i_3025 (.A(in2[11]), .B(in1[31]), .C1(n_2262), .C2(n_1383), 
      .ZN(n_2257));
   OAI211_X1 i_3026 (.A(in2[12]), .B(in1[30]), .C1(n_2259), .C2(n_1384), 
      .ZN(n_2258));
   INV_X1 i_3027 (.A(in2[11]), .ZN(n_2259));
   INV_X1 i_3028 (.A(in2[12]), .ZN(n_2262));
   OAI21_X1 i_3029 (.A(n_2264), .B1(n_2304), .B2(n_2270), .ZN(n_2263));
   NAND2_X1 i_3030 (.A1(n_2305), .A2(n_2266), .ZN(n_2264));
   OAI21_X1 i_3031 (.A(n_2266), .B1(n_2304), .B2(n_2270), .ZN(n_2265));
   NAND2_X1 i_3032 (.A1(n_2304), .A2(n_2270), .ZN(n_2266));
   NOR2_X1 i_3033 (.A1(n_2859), .A2(n_1384), .ZN(n_2270));
   NAND2_X1 i_3034 (.A1(in1[30]), .A2(in2[19]), .ZN(n_2304));
   OAI21_X1 i_3035 (.A(n_2855), .B1(n_2740), .B2(n_2738), .ZN(n_2305));
   NAND2_X1 i_3036 (.A1(in1[29]), .A2(in2[19]), .ZN(n_2738));
   INV_X1 i_3037 (.A(n_2853), .ZN(n_2740));
   OAI211_X1 i_3038 (.A(in2[17]), .B(in1[31]), .C1(n_2859), .C2(n_1383), 
      .ZN(n_2853));
   OAI211_X1 i_3039 (.A(in2[18]), .B(in1[30]), .C1(n_2857), .C2(n_1384), 
      .ZN(n_2855));
   INV_X1 i_3040 (.A(in2[17]), .ZN(n_2857));
   INV_X1 i_3041 (.A(in2[18]), .ZN(n_2859));
   FA_X1 i_3042 (.A(n_735), .B(n_563), .CI(n_562), .CO(n_2863), .S(n_544));
   FA_X1 i_3043 (.A(n_561), .B(n_560), .CI(n_559), .CO(n_546), .S(n_2865));
   FA_X1 i_3044 (.A(n_546), .B(n_558), .CI(n_557), .CO(n_547), .S(n_2893));
   FA_X1 i_3045 (.A(n_555), .B(n_554), .CI(n_553), .CO(n_549), .S(n_2966));
   FA_X1 i_3046 (.A(n_556), .B(n_549), .CI(n_551), .CO(n_2972), .S(n_550));
   FA_X1 i_3047 (.A(n_544), .B(n_547), .CI(n_550), .CO(n_2980), .S(n_2978));
   OAI21_X1 i_3048 (.A(n_2982), .B1(n_3098), .B2(n_3094), .ZN(n_551));
   NAND2_X1 i_3049 (.A1(n_3092), .A2(n_3083), .ZN(n_2982));
   OAI21_X1 i_3050 (.A(n_3205), .B1(n_3203), .B2(n_3193), .ZN(n_553));
   AOI21_X1 i_3051 (.A(n_3207), .B1(n_3208), .B2(n_3206), .ZN(n_554));
   OAI21_X1 i_3052 (.A(n_3287), .B1(n_3213), .B2(n_3212), .ZN(n_555));
   OAI21_X1 i_3053 (.A(n_3292), .B1(n_3291), .B2(n_3289), .ZN(n_556));
   XOR2_X1 i_3054 (.A(n_3099), .B(n_2984), .Z(n_557));
   OAI21_X1 i_3055 (.A(n_3187), .B1(n_3190), .B2(n_3189), .ZN(n_2984));
   XNOR2_X1 i_3056 (.A(n_3084), .B(n_3083), .ZN(n_558));
   OAI21_X1 i_3057 (.A(n_3313), .B1(n_3305), .B2(n_3303), .ZN(n_3083));
   OAI21_X1 i_3058 (.A(n_3092), .B1(n_3098), .B2(n_3094), .ZN(n_3084));
   NAND2_X1 i_3059 (.A1(n_3098), .A2(n_3094), .ZN(n_3092));
   NOR2_X1 i_3060 (.A1(n_3573), .A2(n_1384), .ZN(n_3094));
   NAND2_X1 i_3061 (.A1(in1[30]), .A2(in2[22]), .ZN(n_3098));
   OAI21_X1 i_3062 (.A(n_3401), .B1(n_3392), .B2(n_3390), .ZN(n_559));
   OAI21_X1 i_3063 (.A(n_3488), .B1(n_3486), .B2(n_3402), .ZN(n_560));
   OAI21_X1 i_3064 (.A(n_3566), .B1(n_3565), .B2(n_3562), .ZN(n_561));
   OAI21_X1 i_3065 (.A(n_3569), .B1(n_3568), .B2(n_3567), .ZN(n_562));
   OAI21_X1 i_3066 (.A(n_3187), .B1(n_3100), .B2(n_3099), .ZN(n_563));
   NAND2_X1 i_3067 (.A1(in1[27]), .A2(in2[25]), .ZN(n_3099));
   NOR2_X1 i_3068 (.A1(n_3190), .A2(n_3189), .ZN(n_3100));
   NAND2_X1 i_3069 (.A1(n_3190), .A2(n_3189), .ZN(n_3187));
   AND2_X1 i_3070 (.A1(in1[29]), .A2(in2[23]), .ZN(n_3189));
   NOR2_X1 i_3071 (.A1(n_3574), .A2(n_1580), .ZN(n_3190));
   NAND2_X1 i_3072 (.A1(in1[31]), .A2(in2[22]), .ZN(n_735));
   AND2_X1 i_3073 (.A1(in1[20]), .A2(in2[31]), .ZN(n_3193));
   AOI22_X1 i_3074 (.A1(in1[21]), .A2(in2[30]), .B1(in1[22]), .B2(in2[29]), 
      .ZN(n_3203));
   NAND4_X1 i_3075 (.A1(in1[21]), .A2(in2[30]), .A3(in1[22]), .A4(in2[29]), 
      .ZN(n_3205));
   NAND2_X1 i_3076 (.A1(in1[23]), .A2(in2[28]), .ZN(n_3206));
   AOI22_X1 i_3077 (.A1(in1[24]), .A2(in2[27]), .B1(in1[25]), .B2(in2[26]), 
      .ZN(n_3207));
   NAND4_X1 i_3078 (.A1(in1[25]), .A2(in2[27]), .A3(in1[24]), .A4(in2[26]), 
      .ZN(n_3208));
   NAND2_X1 i_3079 (.A1(in1[26]), .A2(in2[25]), .ZN(n_3212));
   AOI22_X1 i_3080 (.A1(in1[27]), .A2(in2[24]), .B1(in1[28]), .B2(in2[23]), 
      .ZN(n_3213));
   NAND4_X1 i_3081 (.A1(in1[27]), .A2(in2[24]), .A3(in1[28]), .A4(in2[23]), 
      .ZN(n_3287));
   AND2_X1 i_3082 (.A1(in1[21]), .A2(in2[31]), .ZN(n_3289));
   AOI22_X1 i_3083 (.A1(in1[22]), .A2(in2[30]), .B1(in1[23]), .B2(in2[29]), 
      .ZN(n_3291));
   NAND4_X1 i_3084 (.A1(in1[22]), .A2(in2[30]), .A3(in1[23]), .A4(in2[29]), 
      .ZN(n_3292));
   NAND2_X1 i_3085 (.A1(in1[29]), .A2(in2[22]), .ZN(n_3303));
   INV_X1 i_3086 (.A(n_3312), .ZN(n_3305));
   OAI211_X1 i_3087 (.A(in2[20]), .B(in1[31]), .C1(n_3573), .C2(n_1383), 
      .ZN(n_3312));
   OAI211_X1 i_3088 (.A(in2[21]), .B(in1[30]), .C1(n_3572), .C2(n_1384), 
      .ZN(n_3313));
   NAND2_X1 i_3089 (.A1(in1[22]), .A2(in2[28]), .ZN(n_3390));
   AOI22_X1 i_3090 (.A1(in1[23]), .A2(in2[27]), .B1(in1[24]), .B2(in2[26]), 
      .ZN(n_3392));
   NAND4_X1 i_3091 (.A1(in1[23]), .A2(in2[27]), .A3(in1[24]), .A4(in2[26]), 
      .ZN(n_3401));
   NAND2_X1 i_3092 (.A1(in1[25]), .A2(in2[25]), .ZN(n_3402));
   AOI22_X1 i_3093 (.A1(in1[26]), .A2(in2[24]), .B1(in1[27]), .B2(in2[23]), 
      .ZN(n_3486));
   NAND4_X1 i_3094 (.A1(in1[26]), .A2(in2[24]), .A3(in1[27]), .A4(in2[23]), 
      .ZN(n_3488));
   NAND2_X1 i_3095 (.A1(in1[28]), .A2(in2[22]), .ZN(n_3562));
   AOI22_X1 i_3096 (.A1(in1[29]), .A2(in2[21]), .B1(in1[30]), .B2(in2[20]), 
      .ZN(n_3565));
   NAND4_X1 i_3097 (.A1(in1[29]), .A2(in2[21]), .A3(in1[30]), .A4(in2[20]), 
      .ZN(n_3566));
   NAND2_X1 i_3098 (.A1(in1[24]), .A2(in2[28]), .ZN(n_3567));
   AOI22_X1 i_3099 (.A1(in1[25]), .A2(in2[27]), .B1(in1[26]), .B2(in2[26]), 
      .ZN(n_3568));
   NAND4_X1 i_3100 (.A1(in1[25]), .A2(in2[27]), .A3(in1[26]), .A4(in2[26]), 
      .ZN(n_3569));
   INV_X1 i_3101 (.A(in2[20]), .ZN(n_3572));
   INV_X1 i_3102 (.A(in2[21]), .ZN(n_3573));
   INV_X1 i_3103 (.A(in2[24]), .ZN(n_3574));
   OAI21_X1 i_3104 (.A(n_3581), .B1(n_3620), .B2(n_3611), .ZN(n_3579));
   NAND2_X1 i_3105 (.A1(n_3621), .A2(n_3610), .ZN(n_3581));
   OAI21_X1 i_3106 (.A(n_3610), .B1(n_3620), .B2(n_3611), .ZN(n_3607));
   NAND2_X1 i_3107 (.A1(n_3620), .A2(n_3611), .ZN(n_3610));
   NOR2_X1 i_3108 (.A1(n_1384), .A2(n_3574), .ZN(n_3611));
   NAND2_X1 i_3109 (.A1(in1[30]), .A2(in2[25]), .ZN(n_3620));
   OAI21_X1 i_3110 (.A(n_3648), .B1(n_3644), .B2(n_3643), .ZN(n_3621));
   NAND2_X1 i_3111 (.A1(in1[29]), .A2(in2[25]), .ZN(n_3643));
   INV_X1 i_3112 (.A(n_3647), .ZN(n_3644));
   OAI211_X1 i_3113 (.A(in2[23]), .B(in1[31]), .C1(n_1383), .C2(n_3574), 
      .ZN(n_3647));
   OAI211_X1 i_3114 (.A(in2[24]), .B(in1[30]), .C1(n_3649), .C2(n_1384), 
      .ZN(n_3648));
   INV_X1 i_3115 (.A(in2[23]), .ZN(n_3649));
   FA_X1 i_3116 (.A(n_927), .B(n_570), .CI(n_569), .CO(n_3650), .S(n_564));
   FA_X1 i_3117 (.A(n_568), .B(n_567), .CI(n_566), .CO(n_565), .S(n_3651));
   FA_X1 i_3118 (.A(n_571), .B(n_564), .CI(n_565), .CO(n_3655), .S(n_3654));
   XOR2_X1 i_3119 (.A(n_3707), .B(n_3656), .Z(n_566));
   OAI21_X1 i_3120 (.A(n_3709), .B1(n_3729), .B2(n_3710), .ZN(n_3656));
   XNOR2_X1 i_3121 (.A(n_3678), .B(n_3670), .ZN(n_567));
   OAI21_X1 i_3122 (.A(n_3702), .B1(n_3704), .B2(n_3703), .ZN(n_3670));
   OAI21_X1 i_3123 (.A(n_3716), .B1(n_3715), .B2(n_3714), .ZN(n_568));
   OAI22_X1 i_3124 (.A1(n_3704), .A2(n_3703), .B1(n_3701), .B2(n_3677), .ZN(
      n_569));
   INV_X1 i_3125 (.A(n_3678), .ZN(n_3677));
   OAI21_X1 i_3126 (.A(n_3723), .B1(n_3721), .B2(n_3718), .ZN(n_3678));
   INV_X1 i_3127 (.A(n_3702), .ZN(n_3701));
   NAND2_X1 i_3128 (.A1(n_3704), .A2(n_3703), .ZN(n_3702));
   NOR2_X1 i_3129 (.A1(n_3732), .A2(n_1384), .ZN(n_3703));
   NAND2_X1 i_3130 (.A1(in1[30]), .A2(in2[28]), .ZN(n_3704));
   OAI22_X1 i_3131 (.A1(n_3729), .A2(n_3710), .B1(n_3708), .B2(n_3707), .ZN(
      n_570));
   NOR2_X1 i_3132 (.A1(n_1602), .A2(n_1381), .ZN(n_3707));
   INV_X1 i_3133 (.A(n_3709), .ZN(n_3708));
   NAND2_X1 i_3134 (.A1(n_3729), .A2(n_3710), .ZN(n_3709));
   NAND2_X1 i_3135 (.A1(in1[28]), .A2(in2[30]), .ZN(n_3710));
   NAND2_X1 i_3136 (.A1(in1[31]), .A2(in2[28]), .ZN(n_927));
   XNOR2_X1 i_3137 (.A(n_3724), .B(n_3711), .ZN(n_571));
   NOR2_X1 i_3138 (.A1(n_3728), .A2(n_3725), .ZN(n_3711));
   AND2_X1 i_3139 (.A1(in1[26]), .A2(in2[31]), .ZN(n_3714));
   AOI21_X1 i_3140 (.A(n_3717), .B1(in1[28]), .B2(in2[29]), .ZN(n_3715));
   NAND3_X1 i_3141 (.A1(in1[28]), .A2(in2[29]), .A3(n_3717), .ZN(n_3716));
   AND2_X1 i_3142 (.A1(in1[27]), .A2(in2[30]), .ZN(n_3717));
   NAND2_X1 i_3143 (.A1(in1[29]), .A2(in2[28]), .ZN(n_3718));
   INV_X1 i_3144 (.A(n_3722), .ZN(n_3721));
   OAI211_X1 i_3145 (.A(in2[26]), .B(in1[31]), .C1(n_3732), .C2(n_1383), 
      .ZN(n_3722));
   OAI211_X1 i_3146 (.A(in2[27]), .B(in1[30]), .C1(n_3731), .C2(n_1384), 
      .ZN(n_3723));
   NOR2_X1 i_3147 (.A1(n_1602), .A2(n_1580), .ZN(n_3724));
   AOI22_X1 i_3148 (.A1(in1[29]), .A2(in2[30]), .B1(in1[30]), .B2(in2[29]), 
      .ZN(n_3725));
   NOR2_X1 i_3149 (.A1(n_3730), .A2(n_3729), .ZN(n_3728));
   NAND2_X1 i_3150 (.A1(in1[29]), .A2(in2[29]), .ZN(n_3729));
   NAND2_X1 i_3151 (.A1(in1[30]), .A2(in2[30]), .ZN(n_3730));
   INV_X1 i_3152 (.A(in2[26]), .ZN(n_3731));
   INV_X1 i_3153 (.A(in2[27]), .ZN(n_3732));
endmodule

module VerilogMultiplierCircuit(in1, in2, out, ovflag);
   input [31:0]in1;
   input [31:0]in2;
   output [63:0]out;
   output ovflag;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;

   datapath i_0 (.in2(in2), .in1(in1), .out(out));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(ovflag));
   OAI221_X1 i_1_1 (.A(n_1_11), .B1(n_1_6), .B2(n_1_1), .C1(n_1_18), .C2(n_1_13), 
      .ZN(n_1_0));
   NAND4_X1 i_1_2 (.A1(n_1_5), .A2(n_1_4), .A3(n_1_3), .A4(n_1_2), .ZN(n_1_1));
   NOR4_X1 i_1_3 (.A1(in1[18]), .A2(in1[17]), .A3(in1[23]), .A4(in1[20]), 
      .ZN(n_1_2));
   NOR4_X1 i_1_4 (.A1(in1[27]), .A2(in1[24]), .A3(in1[30]), .A4(in1[29]), 
      .ZN(n_1_3));
   NOR4_X1 i_1_5 (.A1(in1[6]), .A2(in1[5]), .A3(in1[3]), .A4(in1[0]), .ZN(n_1_4));
   NOR4_X1 i_1_6 (.A1(in1[10]), .A2(in1[9]), .A3(in1[15]), .A4(in1[12]), 
      .ZN(n_1_5));
   NAND4_X1 i_1_7 (.A1(n_1_10), .A2(n_1_9), .A3(n_1_8), .A4(n_1_7), .ZN(n_1_6));
   NOR4_X1 i_1_8 (.A1(in1[19]), .A2(in1[16]), .A3(in1[22]), .A4(in1[21]), 
      .ZN(n_1_7));
   NOR4_X1 i_1_9 (.A1(in1[26]), .A2(in1[25]), .A3(in1[31]), .A4(in1[28]), 
      .ZN(n_1_8));
   NOR4_X1 i_1_10 (.A1(in1[2]), .A2(in1[1]), .A3(in1[7]), .A4(in1[4]), .ZN(n_1_9));
   NOR4_X1 i_1_11 (.A1(in1[11]), .A2(in1[8]), .A3(in1[14]), .A4(in1[13]), 
      .ZN(n_1_10));
   XOR2_X1 i_1_12 (.A(out[63]), .B(n_1_12), .Z(n_1_11));
   XOR2_X1 i_1_13 (.A(in2[31]), .B(in1[31]), .Z(n_1_12));
   NAND4_X1 i_1_14 (.A1(n_1_17), .A2(n_1_16), .A3(n_1_15), .A4(n_1_14), .ZN(
      n_1_13));
   NOR4_X1 i_1_15 (.A1(in2[7]), .A2(in2[6]), .A3(in2[5]), .A4(in2[4]), .ZN(
      n_1_14));
   NOR4_X1 i_1_16 (.A1(in2[3]), .A2(in2[2]), .A3(in2[1]), .A4(in2[0]), .ZN(
      n_1_15));
   NOR4_X1 i_1_17 (.A1(in2[15]), .A2(in2[14]), .A3(in2[13]), .A4(in2[12]), 
      .ZN(n_1_16));
   NOR4_X1 i_1_18 (.A1(in2[11]), .A2(in2[10]), .A3(in2[9]), .A4(in2[8]), 
      .ZN(n_1_17));
   NAND4_X1 i_1_19 (.A1(n_1_22), .A2(n_1_21), .A3(n_1_20), .A4(n_1_19), .ZN(
      n_1_18));
   NOR4_X1 i_1_20 (.A1(in2[25]), .A2(in2[24]), .A3(in2[27]), .A4(in2[26]), 
      .ZN(n_1_19));
   NOR4_X1 i_1_21 (.A1(in2[29]), .A2(in2[28]), .A3(in2[31]), .A4(in2[30]), 
      .ZN(n_1_20));
   NOR4_X1 i_1_22 (.A1(in2[21]), .A2(in2[20]), .A3(in2[23]), .A4(in2[22]), 
      .ZN(n_1_21));
   NOR4_X1 i_1_23 (.A1(in2[17]), .A2(in2[16]), .A3(in2[19]), .A4(in2[18]), 
      .ZN(n_1_22));
endmodule

module Register__parameterized0(in, clk, out);
   input [63:0]in;
   input clk;
   output [63:0]out;

   DFF_X1 \out_reg[63]  (.D(in[63]), .CK(clk), .Q(out[63]), .QN());
   DFF_X1 \out_reg[62]  (.D(in[62]), .CK(clk), .Q(out[62]), .QN());
   DFF_X1 \out_reg[61]  (.D(in[61]), .CK(clk), .Q(out[61]), .QN());
   DFF_X1 \out_reg[60]  (.D(in[60]), .CK(clk), .Q(out[60]), .QN());
   DFF_X1 \out_reg[59]  (.D(in[59]), .CK(clk), .Q(out[59]), .QN());
   DFF_X1 \out_reg[58]  (.D(in[58]), .CK(clk), .Q(out[58]), .QN());
   DFF_X1 \out_reg[57]  (.D(in[57]), .CK(clk), .Q(out[57]), .QN());
   DFF_X1 \out_reg[56]  (.D(in[56]), .CK(clk), .Q(out[56]), .QN());
   DFF_X1 \out_reg[55]  (.D(in[55]), .CK(clk), .Q(out[55]), .QN());
   DFF_X1 \out_reg[54]  (.D(in[54]), .CK(clk), .Q(out[54]), .QN());
   DFF_X1 \out_reg[53]  (.D(in[53]), .CK(clk), .Q(out[53]), .QN());
   DFF_X1 \out_reg[52]  (.D(in[52]), .CK(clk), .Q(out[52]), .QN());
   DFF_X1 \out_reg[51]  (.D(in[51]), .CK(clk), .Q(out[51]), .QN());
   DFF_X1 \out_reg[50]  (.D(in[50]), .CK(clk), .Q(out[50]), .QN());
   DFF_X1 \out_reg[49]  (.D(in[49]), .CK(clk), .Q(out[49]), .QN());
   DFF_X1 \out_reg[48]  (.D(in[48]), .CK(clk), .Q(out[48]), .QN());
   DFF_X1 \out_reg[47]  (.D(in[47]), .CK(clk), .Q(out[47]), .QN());
   DFF_X1 \out_reg[46]  (.D(in[46]), .CK(clk), .Q(out[46]), .QN());
   DFF_X1 \out_reg[45]  (.D(in[45]), .CK(clk), .Q(out[45]), .QN());
   DFF_X1 \out_reg[44]  (.D(in[44]), .CK(clk), .Q(out[44]), .QN());
   DFF_X1 \out_reg[43]  (.D(in[43]), .CK(clk), .Q(out[43]), .QN());
   DFF_X1 \out_reg[42]  (.D(in[42]), .CK(clk), .Q(out[42]), .QN());
   DFF_X1 \out_reg[41]  (.D(in[41]), .CK(clk), .Q(out[41]), .QN());
   DFF_X1 \out_reg[40]  (.D(in[40]), .CK(clk), .Q(out[40]), .QN());
   DFF_X1 \out_reg[39]  (.D(in[39]), .CK(clk), .Q(out[39]), .QN());
   DFF_X1 \out_reg[38]  (.D(in[38]), .CK(clk), .Q(out[38]), .QN());
   DFF_X1 \out_reg[37]  (.D(in[37]), .CK(clk), .Q(out[37]), .QN());
   DFF_X1 \out_reg[36]  (.D(in[36]), .CK(clk), .Q(out[36]), .QN());
   DFF_X1 \out_reg[35]  (.D(in[35]), .CK(clk), .Q(out[35]), .QN());
   DFF_X1 \out_reg[34]  (.D(in[34]), .CK(clk), .Q(out[34]), .QN());
   DFF_X1 \out_reg[33]  (.D(in[33]), .CK(clk), .Q(out[33]), .QN());
   DFF_X1 \out_reg[32]  (.D(in[32]), .CK(clk), .Q(out[32]), .QN());
   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module VerilogMultiplier(in1, in2, clk, out, ovflag);
   input [31:0]in1;
   input [31:0]in2;
   input clk;
   output [63:0]out;
   output ovflag;

   wire [63:0]result;

   VerilogMultiplierCircuit VerilogMultiplierCircuitInst (.in1(in1), .in2(in2), 
      .out(result), .ovflag(ovflag));
   Register__parameterized0 Register_inst3 (.in(result), .clk(clk), .out(out));
endmodule
