/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Mon Oct 31 16:36:24 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1885500826 */

module FA__0_5(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_9(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_13(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_17(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_21(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_25(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_29(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_33(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_37(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_41(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_45(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_49(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_53(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_57(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_61(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_65(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_69(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_73(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_77(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_81(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_85(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_89(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_93(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_97(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_101(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_105(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_109(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_113(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_117(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_121(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_125(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA(in1, in2, sum, cout);
   input [31:0]in1;
   input [31:0]in2;
   output [31:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;

   FA__0_5 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(n_0_0));
   FA__0_9 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(n_0_0), 
      .sum(sum[1]), .cout(n_0_1));
   FA__0_13 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(n_0_1), 
      .sum(sum[2]), .cout(n_0_2));
   FA__0_17 genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(n_0_2), 
      .sum(sum[3]), .cout(n_0_3));
   FA__0_21 genblk1_4_full_adder_inst (.in1(in1[4]), .in2(in2[4]), .cin(n_0_3), 
      .sum(sum[4]), .cout(n_0_4));
   FA__0_25 genblk1_5_full_adder_inst (.in1(in1[5]), .in2(in2[5]), .cin(n_0_4), 
      .sum(sum[5]), .cout(n_0_5));
   FA__0_29 genblk1_6_full_adder_inst (.in1(in1[6]), .in2(in2[6]), .cin(n_0_5), 
      .sum(sum[6]), .cout(n_0_6));
   FA__0_33 genblk1_7_full_adder_inst (.in1(in1[7]), .in2(in2[7]), .cin(n_0_6), 
      .sum(sum[7]), .cout(n_0_7));
   FA__0_37 genblk1_8_full_adder_inst (.in1(in1[8]), .in2(in2[8]), .cin(n_0_7), 
      .sum(sum[8]), .cout(n_0_8));
   FA__0_41 genblk1_9_full_adder_inst (.in1(in1[9]), .in2(in2[9]), .cin(n_0_8), 
      .sum(sum[9]), .cout(n_0_9));
   FA__0_45 genblk1_10_full_adder_inst (.in1(in1[10]), .in2(in2[10]), .cin(n_0_9), 
      .sum(sum[10]), .cout(n_0_10));
   FA__0_49 genblk1_11_full_adder_inst (.in1(in1[11]), .in2(in2[11]), .cin(
      n_0_10), .sum(sum[11]), .cout(n_0_11));
   FA__0_53 genblk1_12_full_adder_inst (.in1(in1[12]), .in2(in2[12]), .cin(
      n_0_11), .sum(sum[12]), .cout(n_0_12));
   FA__0_57 genblk1_13_full_adder_inst (.in1(in1[13]), .in2(in2[13]), .cin(
      n_0_12), .sum(sum[13]), .cout(n_0_13));
   FA__0_61 genblk1_14_full_adder_inst (.in1(in1[14]), .in2(in2[14]), .cin(
      n_0_13), .sum(sum[14]), .cout(n_0_14));
   FA__0_65 genblk1_15_full_adder_inst (.in1(in1[15]), .in2(in2[15]), .cin(
      n_0_14), .sum(sum[15]), .cout(n_0_15));
   FA__0_69 genblk1_16_full_adder_inst (.in1(in1[16]), .in2(in2[16]), .cin(
      n_0_15), .sum(sum[16]), .cout(n_0_16));
   FA__0_73 genblk1_17_full_adder_inst (.in1(in1[17]), .in2(in2[17]), .cin(
      n_0_16), .sum(sum[17]), .cout(n_0_17));
   FA__0_77 genblk1_18_full_adder_inst (.in1(in1[18]), .in2(in2[18]), .cin(
      n_0_17), .sum(sum[18]), .cout(n_0_18));
   FA__0_81 genblk1_19_full_adder_inst (.in1(in1[19]), .in2(in2[19]), .cin(
      n_0_18), .sum(sum[19]), .cout(n_0_19));
   FA__0_85 genblk1_20_full_adder_inst (.in1(in1[20]), .in2(in2[20]), .cin(
      n_0_19), .sum(sum[20]), .cout(n_0_20));
   FA__0_89 genblk1_21_full_adder_inst (.in1(in1[21]), .in2(in2[21]), .cin(
      n_0_20), .sum(sum[21]), .cout(n_0_21));
   FA__0_93 genblk1_22_full_adder_inst (.in1(in1[22]), .in2(in2[22]), .cin(
      n_0_21), .sum(sum[22]), .cout(n_0_22));
   FA__0_97 genblk1_23_full_adder_inst (.in1(in1[23]), .in2(in2[23]), .cin(
      n_0_22), .sum(sum[23]), .cout(n_0_23));
   FA__0_101 genblk1_24_full_adder_inst (.in1(in1[24]), .in2(in2[24]), .cin(
      n_0_23), .sum(sum[24]), .cout(n_0_24));
   FA__0_105 genblk1_25_full_adder_inst (.in1(in1[25]), .in2(in2[25]), .cin(
      n_0_24), .sum(sum[25]), .cout(n_0_25));
   FA__0_109 genblk1_26_full_adder_inst (.in1(in1[26]), .in2(in2[26]), .cin(
      n_0_25), .sum(sum[26]), .cout(n_0_26));
   FA__0_113 genblk1_27_full_adder_inst (.in1(in1[27]), .in2(in2[27]), .cin(
      n_0_26), .sum(sum[27]), .cout(n_0_27));
   FA__0_117 genblk1_28_full_adder_inst (.in1(in1[28]), .in2(in2[28]), .cin(
      n_0_27), .sum(sum[28]), .cout(n_0_28));
   FA__0_121 genblk1_29_full_adder_inst (.in1(in1[29]), .in2(in2[29]), .cin(
      n_0_28), .sum(sum[29]), .cout(n_0_29));
   FA__0_125 genblk1_30_full_adder_inst (.in1(in1[30]), .in2(in2[30]), .cin(
      n_0_29), .sum(sum[30]), .cout(n_0_30));
   FA genblk1_31_full_adder_inst (.in1(in1[31]), .in2(in2[31]), .cin(n_0_30), 
      .sum(sum[31]), .cout(cout));
endmodule
