module LZeros(input[23:0]in,output[4:0]out);
assign out=(in[23]==1)?5'b0:
(in[22]==1)?5'b00001:
(in[21]==1)?5'b00010:
(in[20]==1)?5'b00011:
(in[19]==1)?5'b00100:
(in[18]==1)?5'b00101:
(in[17]==1)?5'b00110:
(in[16]==1)?5'b00111:
(in[15]==1)?5'b01000:
(in[14]==1)?5'b01001:
(in[13]==1)?5'b01010:
(in[12]==1)?5'b01011:
(in[11]==1)?5'b01100:
(in[10]==1)?5'b01101:
(in[9]==1)?5'b01110:
(in[8]==1)?5'b01111:
(in[7]==1)?5'b10000:
(in[6]==1)?5'b10001:
(in[5]==1)?5'b10010:
(in[4]==1)?5'b10011:
(in[3]==1)?5'b10100:
(in[2]==1)?5'b10101:
(in[1]==1)?5'b10110:
(in[0]==1)?5'b10111:5'b0;
endmodule
