
// 	Thu Dec 22 04:27:06 2022
//	vlsi
//	localhost.localdomain

module Register__parameterized0 (clk_CTSPP_157, clk_CTSPP_154, clk_CTSPP_156, clk_CTSPP_159, 
    in, clk, out);

output [63:0] out;
output clk_CTSPP_157;
input clk;
input [63:0] in;
input clk_CTSPP_154;
input clk_CTSPP_156;
input clk_CTSPP_159;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk_CTSPP_156), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk_CTSPP_156), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk_CTSPP_156), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk_CTSPP_156), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk_CTSPP_156), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk_CTSPP_157), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk_CTSPP_157), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk_CTSPP_157), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk_CTSPP_157), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk_CTSPP_157), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk_CTSPP_157), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk_CTSPP_157), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk_CTSPP_157), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk_CTSPP_157), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk_CTSPP_157), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk_CTSPP_157), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk_CTSPP_157), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk_CTSPP_157), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk_CTSPP_156), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk_CTSPP_156), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk_CTSPP_156), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk_CTSPP_156), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk_CTSPP_156), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk_CTSPP_156), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk_CTSPP_156), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk_CTSPP_156), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk_CTSPP_156), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk_CTSPP_156), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk_CTSPP_156), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk_CTSPP_156), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk_CTSPP_157), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk_CTSPP_157), .D (in[31]));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (clk_CTSPP_157), .D (in[32]));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (clk_CTSPP_157), .D (in[33]));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (clk_CTSPP_157), .D (in[34]));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (clk_CTSPP_157), .D (in[35]));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (clk_CTSPP_157), .D (in[36]));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (clk_CTSPP_157), .D (in[37]));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (clk_CTSPP_157), .D (in[38]));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (clk_CTSPP_157), .D (in[39]));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (clk_CTSPP_157), .D (in[40]));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (clk_CTSPP_157), .D (in[41]));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (clk_CTSPP_157), .D (in[42]));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (clk_CTSPP_157), .D (in[43]));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (clk_CTSPP_157), .D (in[44]));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (clk_CTSPP_157), .D (in[45]));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (clk_CTSPP_154), .D (in[46]));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (clk_CTSPP_157), .D (in[47]));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (clk_CTSPP_154), .D (in[48]));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (clk_CTSPP_154), .D (in[49]));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (clk_CTSPP_154), .D (in[50]));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (clk_CTSPP_154), .D (in[51]));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (clk_CTSPP_154), .D (in[52]));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (clk_CTSPP_154), .D (in[53]));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (clk_CTSPP_154), .D (in[54]));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (clk_CTSPP_154), .D (in[55]));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (clk_CTSPP_154), .D (in[56]));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (clk_CTSPP_154), .D (in[57]));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (clk_CTSPP_154), .D (in[58]));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (clk_CTSPP_154), .D (in[59]));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (clk_CTSPP_154), .D (in[60]));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (clk_CTSPP_154), .D (in[61]));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (clk_CTSPP_154), .D (in[62]));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (clk_CTSPP_154), .D (in[63]));
CLKBUF_X3 CTS_L2_c25 (.Z (clk_CTSPP_157), .A (clk_CTSPP_159));

endmodule //Register__parameterized0

module datapath__0_10 (p_0, acc_out, acc_out1);

output [63:0] acc_out1;
input [63:0] acc_out;
input [63:0] p_0;
wire n_0;
wire n_366;
wire n_1;
wire n_365;
wire n_364;
wire n_2;
wire n_369;
wire n_363;
wire n_3;
wire n_370;
wire n_376;
wire n_372;
wire n_361;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_358;
wire n_349;
wire n_11;
wire n_5;
wire n_359;
wire n_353;
wire n_8;
wire n_356;
wire n_354;
wire n_360;
wire n_351;
wire n_347;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_344;
wire n_335;
wire n_19;
wire n_13;
wire n_345;
wire n_339;
wire n_16;
wire n_342;
wire n_340;
wire n_346;
wire n_337;
wire n_333;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_330;
wire n_321;
wire n_27;
wire n_21;
wire n_331;
wire n_325;
wire n_24;
wire n_328;
wire n_326;
wire n_332;
wire n_323;
wire n_319;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_285;
wire n_275;
wire n_35;
wire n_29;
wire n_284;
wire n_287;
wire n_277;
wire n_32;
wire n_286;
wire n_282;
wire n_279;
wire n_289;
wire n_63;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_313;
wire n_257;
wire n_43;
wire n_37;
wire n_312;
wire n_315;
wire n_259;
wire n_40;
wire n_314;
wire n_318;
wire n_261;
wire n_317;
wire n_61;
wire n_50;
wire n_49;
wire n_46;
wire n_47;
wire n_44;
wire n_296;
wire n_269;
wire n_51;
wire n_45;
wire n_295;
wire n_298;
wire n_271;
wire n_48;
wire n_297;
wire n_293;
wire n_273;
wire n_300;
wire n_59;
wire n_58;
wire n_57;
wire n_54;
wire n_55;
wire n_52;
wire n_305;
wire n_263;
wire n_65;
wire n_53;
wire n_304;
wire n_307;
wire n_266;
wire n_56;
wire n_306;
wire n_302;
wire n_267;
wire n_60;
wire n_268;
wire n_292;
wire n_62;
wire n_256;
wire n_310;
wire n_64;
wire n_274;
wire n_281;
wire n_308;
wire n_377;
wire n_373;
wire n_254;
wire n_72;
wire n_71;
wire n_68;
wire n_69;
wire n_66;
wire n_223;
wire n_213;
wire n_73;
wire n_67;
wire n_222;
wire n_225;
wire n_215;
wire n_70;
wire n_224;
wire n_220;
wire n_217;
wire n_227;
wire n_101;
wire n_80;
wire n_79;
wire n_76;
wire n_77;
wire n_74;
wire n_248;
wire n_206;
wire n_81;
wire n_75;
wire n_247;
wire n_250;
wire n_208;
wire n_78;
wire n_249;
wire n_253;
wire n_210;
wire n_252;
wire n_99;
wire n_88;
wire n_87;
wire n_84;
wire n_85;
wire n_82;
wire n_234;
wire n_192;
wire n_89;
wire n_83;
wire n_233;
wire n_236;
wire n_194;
wire n_86;
wire n_235;
wire n_231;
wire n_196;
wire n_238;
wire n_98;
wire n_97;
wire n_95;
wire n_94;
wire n_91;
wire n_90;
wire n_202;
wire n_242;
wire n_199;
wire n_103;
wire n_92;
wire n_93;
wire n_241;
wire n_200;
wire n_96;
wire n_243;
wire n_203;
wire n_204;
wire n_191;
wire n_230;
wire n_100;
wire n_205;
wire n_245;
wire n_102;
wire n_212;
wire n_219;
wire n_244;
wire n_189;
wire n_110;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_186;
wire n_177;
wire n_111;
wire n_105;
wire n_187;
wire n_181;
wire n_108;
wire n_184;
wire n_182;
wire n_188;
wire n_179;
wire n_175;
wire n_118;
wire n_117;
wire n_114;
wire n_115;
wire n_112;
wire n_164;
wire n_154;
wire n_119;
wire n_113;
wire n_163;
wire n_166;
wire n_156;
wire n_116;
wire n_165;
wire n_161;
wire n_158;
wire n_168;
wire n_128;
wire n_127;
wire n_125;
wire n_124;
wire n_121;
wire n_120;
wire n_149;
wire n_172;
wire n_145;
wire n_129;
wire n_122;
wire n_123;
wire n_171;
wire n_146;
wire n_126;
wire n_173;
wire n_150;
wire n_151;
wire n_153;
wire n_160;
wire n_174;
wire n_143;
wire n_142;
wire n_140;
wire n_136;
wire n_141;
wire n_135;
wire n_131;
wire n_130;
wire n_137;
wire n_139;
wire n_133;
wire n_132;
wire n_134;
wire n_138;
wire n_379;
wire n_375;
wire n_371;
wire n_147;
wire n_144;
wire n_152;
wire n_159;
wire n_378;
wire n_374;
wire n_148;
wire n_170;
wire n_169;
wire n_155;
wire n_167;
wire n_162;
wire n_157;
wire n_176;
wire n_180;
wire n_183;
wire n_178;
wire n_185;
wire n_211;
wire n_190;
wire n_218;
wire n_197;
wire n_239;
wire n_229;
wire n_193;
wire n_237;
wire n_232;
wire n_195;
wire n_198;
wire n_201;
wire n_240;
wire n_207;
wire n_251;
wire n_246;
wire n_209;
wire n_228;
wire n_214;
wire n_226;
wire n_221;
wire n_216;
wire n_262;
wire n_255;
wire n_280;
wire n_290;
wire n_291;
wire n_301;
wire n_258;
wire n_316;
wire n_311;
wire n_260;
wire n_303;
wire n_265;
wire n_309;
wire n_264;
wire n_270;
wire n_299;
wire n_294;
wire n_272;
wire n_276;
wire n_288;
wire n_283;
wire n_278;
wire n_320;
wire n_324;
wire n_327;
wire n_322;
wire n_329;
wire n_334;
wire n_338;
wire n_341;
wire n_336;
wire n_343;
wire n_348;
wire n_352;
wire n_355;
wire n_350;
wire n_357;
wire n_362;
wire n_368;
wire n_367;


INV_X1 i_443 (.ZN (n_379), .A (p_0[61]));
INV_X1 i_442 (.ZN (n_378), .A (p_0[59]));
INV_X1 i_441 (.ZN (n_377), .A (p_0[31]));
INV_X1 i_440 (.ZN (n_376), .A (p_0[3]));
INV_X1 i_439 (.ZN (n_375), .A (acc_out[61]));
INV_X1 i_438 (.ZN (n_374), .A (acc_out[59]));
INV_X1 i_437 (.ZN (n_373), .A (acc_out[31]));
INV_X1 i_436 (.ZN (n_372), .A (acc_out[3]));
NOR2_X1 i_435 (.ZN (n_371), .A1 (p_0[60]), .A2 (acc_out[60]));
NAND2_X1 i_434 (.ZN (n_370), .A1 (n_376), .A2 (n_372));
NAND2_X1 i_433 (.ZN (n_369), .A1 (p_0[2]), .A2 (acc_out[2]));
INV_X1 i_432 (.ZN (n_368), .A (n_369));
NOR2_X1 i_431 (.ZN (n_367), .A1 (p_0[1]), .A2 (acc_out[1]));
NAND2_X1 i_430 (.ZN (n_366), .A1 (p_0[0]), .A2 (acc_out[0]));
NAND2_X1 i_429 (.ZN (n_365), .A1 (p_0[1]), .A2 (acc_out[1]));
AOI21_X1 i_428 (.ZN (n_364), .A (n_367), .B1 (n_366), .B2 (n_365));
OAI22_X1 i_427 (.ZN (n_363), .A1 (p_0[2]), .A2 (acc_out[2]), .B1 (n_368), .B2 (n_364));
OAI21_X1 i_426 (.ZN (n_362), .A (n_363), .B1 (n_376), .B2 (n_372));
NAND2_X1 i_425 (.ZN (n_361), .A1 (n_370), .A2 (n_362));
NOR2_X1 i_424 (.ZN (n_360), .A1 (p_0[7]), .A2 (acc_out[7]));
NOR2_X1 i_423 (.ZN (n_359), .A1 (p_0[5]), .A2 (acc_out[5]));
NOR2_X1 i_422 (.ZN (n_358), .A1 (p_0[6]), .A2 (acc_out[6]));
OR3_X1 i_421 (.ZN (n_357), .A1 (n_360), .A2 (n_358), .A3 (n_359));
NOR2_X1 i_420 (.ZN (n_356), .A1 (p_0[4]), .A2 (acc_out[4]));
NOR3_X1 i_419 (.ZN (n_355), .A1 (n_357), .A2 (n_356), .A3 (n_361));
NAND2_X1 i_418 (.ZN (n_354), .A1 (p_0[4]), .A2 (acc_out[4]));
NAND2_X1 i_417 (.ZN (n_353), .A1 (p_0[5]), .A2 (acc_out[5]));
AOI21_X1 i_416 (.ZN (n_352), .A (n_357), .B1 (n_354), .B2 (n_353));
AND2_X1 i_415 (.ZN (n_351), .A1 (p_0[7]), .A2 (acc_out[7]));
NAND2_X1 i_414 (.ZN (n_350), .A1 (p_0[6]), .A2 (acc_out[6]));
INV_X1 i_413 (.ZN (n_349), .A (n_350));
NOR2_X1 i_412 (.ZN (n_348), .A1 (n_360), .A2 (n_350));
NOR4_X1 i_411 (.ZN (n_347), .A1 (n_351), .A2 (n_348), .A3 (n_352), .A4 (n_355));
NOR2_X1 i_410 (.ZN (n_346), .A1 (p_0[11]), .A2 (acc_out[11]));
NOR2_X1 i_409 (.ZN (n_345), .A1 (p_0[9]), .A2 (acc_out[9]));
NOR2_X1 i_408 (.ZN (n_344), .A1 (p_0[10]), .A2 (acc_out[10]));
OR3_X1 i_407 (.ZN (n_343), .A1 (n_346), .A2 (n_344), .A3 (n_345));
NOR2_X1 i_406 (.ZN (n_342), .A1 (p_0[8]), .A2 (acc_out[8]));
NOR3_X1 i_405 (.ZN (n_341), .A1 (n_343), .A2 (n_342), .A3 (n_347));
NAND2_X1 i_404 (.ZN (n_340), .A1 (p_0[8]), .A2 (acc_out[8]));
NAND2_X1 i_403 (.ZN (n_339), .A1 (p_0[9]), .A2 (acc_out[9]));
AOI21_X1 i_402 (.ZN (n_338), .A (n_343), .B1 (n_340), .B2 (n_339));
AND2_X1 i_401 (.ZN (n_337), .A1 (p_0[11]), .A2 (acc_out[11]));
NAND2_X1 i_400 (.ZN (n_336), .A1 (p_0[10]), .A2 (acc_out[10]));
INV_X1 i_399 (.ZN (n_335), .A (n_336));
NOR2_X1 i_398 (.ZN (n_334), .A1 (n_346), .A2 (n_336));
NOR4_X1 i_397 (.ZN (n_333), .A1 (n_337), .A2 (n_334), .A3 (n_338), .A4 (n_341));
NOR2_X1 i_396 (.ZN (n_332), .A1 (p_0[15]), .A2 (acc_out[15]));
NOR2_X1 i_395 (.ZN (n_331), .A1 (p_0[13]), .A2 (acc_out[13]));
NOR2_X1 i_394 (.ZN (n_330), .A1 (p_0[14]), .A2 (acc_out[14]));
OR3_X1 i_393 (.ZN (n_329), .A1 (n_332), .A2 (n_330), .A3 (n_331));
NOR2_X1 i_392 (.ZN (n_328), .A1 (p_0[12]), .A2 (acc_out[12]));
NOR3_X1 i_391 (.ZN (n_327), .A1 (n_329), .A2 (n_328), .A3 (n_333));
NAND2_X1 i_390 (.ZN (n_326), .A1 (p_0[12]), .A2 (acc_out[12]));
NAND2_X1 i_389 (.ZN (n_325), .A1 (p_0[13]), .A2 (acc_out[13]));
AOI21_X1 i_388 (.ZN (n_324), .A (n_329), .B1 (n_326), .B2 (n_325));
AND2_X1 i_387 (.ZN (n_323), .A1 (p_0[15]), .A2 (acc_out[15]));
NAND2_X1 i_386 (.ZN (n_322), .A1 (p_0[14]), .A2 (acc_out[14]));
INV_X1 i_385 (.ZN (n_321), .A (n_322));
NOR2_X1 i_384 (.ZN (n_320), .A1 (n_332), .A2 (n_322));
NOR4_X1 i_383 (.ZN (n_319), .A1 (n_323), .A2 (n_320), .A3 (n_324), .A4 (n_327));
NOR2_X1 i_382 (.ZN (n_318), .A1 (p_0[20]), .A2 (acc_out[20]));
NOR2_X1 i_381 (.ZN (n_317), .A1 (p_0[23]), .A2 (acc_out[23]));
INV_X1 i_380 (.ZN (n_316), .A (n_317));
NOR2_X1 i_379 (.ZN (n_315), .A1 (p_0[21]), .A2 (acc_out[21]));
INV_X1 i_378 (.ZN (n_314), .A (n_315));
NOR2_X1 i_377 (.ZN (n_313), .A1 (p_0[22]), .A2 (acc_out[22]));
INV_X1 i_376 (.ZN (n_312), .A (n_313));
NAND3_X1 i_375 (.ZN (n_311), .A1 (n_316), .A2 (n_312), .A3 (n_314));
OR2_X1 i_374 (.ZN (n_310), .A1 (n_318), .A2 (n_311));
NOR2_X1 i_373 (.ZN (n_309), .A1 (p_0[31]), .A2 (acc_out[31]));
INV_X1 i_372 (.ZN (n_308), .A (n_309));
NOR2_X1 i_371 (.ZN (n_307), .A1 (p_0[29]), .A2 (acc_out[29]));
INV_X1 i_370 (.ZN (n_306), .A (n_307));
NOR2_X1 i_369 (.ZN (n_305), .A1 (p_0[30]), .A2 (acc_out[30]));
INV_X1 i_368 (.ZN (n_304), .A (n_305));
NAND3_X1 i_367 (.ZN (n_303), .A1 (n_308), .A2 (n_304), .A3 (n_306));
NOR2_X1 i_366 (.ZN (n_302), .A1 (p_0[28]), .A2 (acc_out[28]));
OR2_X1 i_365 (.ZN (n_301), .A1 (n_303), .A2 (n_302));
NOR2_X1 i_364 (.ZN (n_300), .A1 (p_0[27]), .A2 (acc_out[27]));
INV_X1 i_363 (.ZN (n_299), .A (n_300));
NOR2_X1 i_362 (.ZN (n_298), .A1 (p_0[25]), .A2 (acc_out[25]));
INV_X1 i_361 (.ZN (n_297), .A (n_298));
NOR2_X1 i_360 (.ZN (n_296), .A1 (p_0[26]), .A2 (acc_out[26]));
INV_X1 i_359 (.ZN (n_295), .A (n_296));
NAND3_X1 i_358 (.ZN (n_294), .A1 (n_299), .A2 (n_295), .A3 (n_297));
NOR2_X1 i_357 (.ZN (n_293), .A1 (p_0[24]), .A2 (acc_out[24]));
OR2_X1 i_356 (.ZN (n_292), .A1 (n_294), .A2 (n_293));
OR2_X1 i_355 (.ZN (n_291), .A1 (n_301), .A2 (n_292));
OR2_X1 i_354 (.ZN (n_290), .A1 (n_310), .A2 (n_291));
NOR2_X1 i_353 (.ZN (n_289), .A1 (p_0[19]), .A2 (acc_out[19]));
INV_X1 i_352 (.ZN (n_288), .A (n_289));
NOR2_X1 i_351 (.ZN (n_287), .A1 (p_0[17]), .A2 (acc_out[17]));
INV_X1 i_350 (.ZN (n_286), .A (n_287));
NOR2_X1 i_349 (.ZN (n_285), .A1 (p_0[18]), .A2 (acc_out[18]));
INV_X1 i_348 (.ZN (n_284), .A (n_285));
NAND3_X1 i_347 (.ZN (n_283), .A1 (n_288), .A2 (n_284), .A3 (n_286));
NOR2_X1 i_346 (.ZN (n_282), .A1 (p_0[16]), .A2 (acc_out[16]));
OR2_X1 i_345 (.ZN (n_281), .A1 (n_283), .A2 (n_282));
NOR3_X1 i_344 (.ZN (n_280), .A1 (n_290), .A2 (n_281), .A3 (n_319));
NAND2_X1 i_343 (.ZN (n_279), .A1 (p_0[16]), .A2 (acc_out[16]));
NAND2_X1 i_342 (.ZN (n_278), .A1 (p_0[17]), .A2 (acc_out[17]));
INV_X1 i_341 (.ZN (n_277), .A (n_278));
AOI21_X1 i_340 (.ZN (n_276), .A (n_283), .B1 (n_279), .B2 (n_278));
AND2_X1 i_339 (.ZN (n_275), .A1 (p_0[18]), .A2 (acc_out[18]));
AOI221_X1 i_338 (.ZN (n_274), .A (n_276), .B1 (p_0[19]), .B2 (acc_out[19]), .C1 (n_288), .C2 (n_275));
NAND2_X1 i_337 (.ZN (n_273), .A1 (p_0[24]), .A2 (acc_out[24]));
NAND2_X1 i_336 (.ZN (n_272), .A1 (p_0[25]), .A2 (acc_out[25]));
INV_X1 i_335 (.ZN (n_271), .A (n_272));
AOI21_X1 i_334 (.ZN (n_270), .A (n_294), .B1 (n_273), .B2 (n_272));
AND2_X1 i_333 (.ZN (n_269), .A1 (p_0[26]), .A2 (acc_out[26]));
AOI221_X1 i_332 (.ZN (n_268), .A (n_270), .B1 (p_0[27]), .B2 (acc_out[27]), .C1 (n_299), .C2 (n_269));
NAND2_X1 i_331 (.ZN (n_267), .A1 (p_0[28]), .A2 (acc_out[28]));
AND2_X1 i_330 (.ZN (n_266), .A1 (p_0[29]), .A2 (acc_out[29]));
AOI21_X1 i_329 (.ZN (n_265), .A (n_266), .B1 (p_0[28]), .B2 (acc_out[28]));
NAND2_X1 i_328 (.ZN (n_264), .A1 (p_0[30]), .A2 (acc_out[30]));
INV_X1 i_327 (.ZN (n_263), .A (n_264));
OAI222_X1 i_326 (.ZN (n_262), .A1 (n_303), .A2 (n_265), .B1 (n_309), .B2 (n_264), .C1 (n_377), .C2 (n_373));
NAND2_X1 i_325 (.ZN (n_261), .A1 (p_0[20]), .A2 (acc_out[20]));
NAND2_X1 i_324 (.ZN (n_260), .A1 (p_0[21]), .A2 (acc_out[21]));
INV_X1 i_323 (.ZN (n_259), .A (n_260));
AOI21_X1 i_322 (.ZN (n_258), .A (n_311), .B1 (n_261), .B2 (n_260));
AND2_X1 i_321 (.ZN (n_257), .A1 (p_0[22]), .A2 (acc_out[22]));
AOI221_X1 i_320 (.ZN (n_256), .A (n_258), .B1 (p_0[23]), .B2 (acc_out[23]), .C1 (n_316), .C2 (n_257));
OAI222_X1 i_319 (.ZN (n_255), .A1 (n_290), .A2 (n_274), .B1 (n_291), .B2 (n_256), .C1 (n_301), .C2 (n_268));
NOR3_X1 i_318 (.ZN (n_254), .A1 (n_262), .A2 (n_255), .A3 (n_280));
NOR2_X1 i_317 (.ZN (n_253), .A1 (p_0[36]), .A2 (acc_out[36]));
NOR2_X1 i_316 (.ZN (n_252), .A1 (p_0[39]), .A2 (acc_out[39]));
INV_X1 i_315 (.ZN (n_251), .A (n_252));
NOR2_X1 i_314 (.ZN (n_250), .A1 (p_0[37]), .A2 (acc_out[37]));
INV_X1 i_313 (.ZN (n_249), .A (n_250));
NOR2_X1 i_312 (.ZN (n_248), .A1 (p_0[38]), .A2 (acc_out[38]));
INV_X1 i_311 (.ZN (n_247), .A (n_248));
NAND3_X1 i_310 (.ZN (n_246), .A1 (n_251), .A2 (n_247), .A3 (n_249));
OR2_X1 i_309 (.ZN (n_245), .A1 (n_253), .A2 (n_246));
NOR2_X1 i_308 (.ZN (n_244), .A1 (p_0[47]), .A2 (acc_out[47]));
NOR2_X1 i_307 (.ZN (n_243), .A1 (p_0[45]), .A2 (acc_out[45]));
NOR2_X1 i_306 (.ZN (n_242), .A1 (p_0[46]), .A2 (acc_out[46]));
NOR2_X1 i_305 (.ZN (n_241), .A1 (n_243), .A2 (n_242));
NOR3_X1 i_304 (.ZN (n_240), .A1 (n_244), .A2 (n_242), .A3 (n_243));
OAI21_X1 i_303 (.ZN (n_239), .A (n_240), .B1 (p_0[44]), .B2 (acc_out[44]));
NOR2_X1 i_302 (.ZN (n_238), .A1 (p_0[43]), .A2 (acc_out[43]));
INV_X1 i_301 (.ZN (n_237), .A (n_238));
NOR2_X1 i_300 (.ZN (n_236), .A1 (p_0[41]), .A2 (acc_out[41]));
INV_X1 i_299 (.ZN (n_235), .A (n_236));
NOR2_X1 i_298 (.ZN (n_234), .A1 (p_0[42]), .A2 (acc_out[42]));
INV_X1 i_297 (.ZN (n_233), .A (n_234));
NAND3_X1 i_296 (.ZN (n_232), .A1 (n_237), .A2 (n_233), .A3 (n_235));
NOR2_X1 i_295 (.ZN (n_231), .A1 (p_0[40]), .A2 (acc_out[40]));
OR2_X1 i_294 (.ZN (n_230), .A1 (n_232), .A2 (n_231));
OR2_X1 i_293 (.ZN (n_229), .A1 (n_239), .A2 (n_230));
OR2_X1 i_292 (.ZN (n_228), .A1 (n_245), .A2 (n_229));
NOR2_X1 i_291 (.ZN (n_227), .A1 (p_0[35]), .A2 (acc_out[35]));
INV_X1 i_290 (.ZN (n_226), .A (n_227));
NOR2_X1 i_289 (.ZN (n_225), .A1 (p_0[33]), .A2 (acc_out[33]));
INV_X1 i_288 (.ZN (n_224), .A (n_225));
NOR2_X1 i_287 (.ZN (n_223), .A1 (p_0[34]), .A2 (acc_out[34]));
INV_X1 i_286 (.ZN (n_222), .A (n_223));
NAND3_X1 i_285 (.ZN (n_221), .A1 (n_226), .A2 (n_222), .A3 (n_224));
NOR2_X1 i_284 (.ZN (n_220), .A1 (p_0[32]), .A2 (acc_out[32]));
OR2_X1 i_283 (.ZN (n_219), .A1 (n_221), .A2 (n_220));
NOR3_X1 i_282 (.ZN (n_218), .A1 (n_228), .A2 (n_219), .A3 (n_254));
NAND2_X1 i_281 (.ZN (n_217), .A1 (p_0[32]), .A2 (acc_out[32]));
NAND2_X1 i_280 (.ZN (n_216), .A1 (p_0[33]), .A2 (acc_out[33]));
INV_X1 i_279 (.ZN (n_215), .A (n_216));
AOI21_X1 i_278 (.ZN (n_214), .A (n_221), .B1 (n_217), .B2 (n_216));
AND2_X1 i_277 (.ZN (n_213), .A1 (p_0[34]), .A2 (acc_out[34]));
AOI221_X1 i_276 (.ZN (n_212), .A (n_214), .B1 (p_0[35]), .B2 (acc_out[35]), .C1 (n_226), .C2 (n_213));
NOR2_X1 i_275 (.ZN (n_211), .A1 (n_228), .A2 (n_212));
NAND2_X1 i_274 (.ZN (n_210), .A1 (p_0[36]), .A2 (acc_out[36]));
NAND2_X1 i_273 (.ZN (n_209), .A1 (p_0[37]), .A2 (acc_out[37]));
INV_X1 i_272 (.ZN (n_208), .A (n_209));
AOI21_X1 i_271 (.ZN (n_207), .A (n_246), .B1 (n_210), .B2 (n_209));
AND2_X1 i_270 (.ZN (n_206), .A1 (p_0[38]), .A2 (acc_out[38]));
AOI221_X1 i_269 (.ZN (n_205), .A (n_207), .B1 (p_0[39]), .B2 (acc_out[39]), .C1 (n_251), .C2 (n_206));
NAND2_X1 i_268 (.ZN (n_204), .A1 (p_0[44]), .A2 (acc_out[44]));
INV_X1 i_267 (.ZN (n_203), .A (n_204));
AND2_X1 i_266 (.ZN (n_202), .A1 (p_0[45]), .A2 (acc_out[45]));
OAI21_X1 i_265 (.ZN (n_201), .A (n_240), .B1 (n_203), .B2 (n_202));
NAND2_X1 i_264 (.ZN (n_200), .A1 (p_0[46]), .A2 (acc_out[46]));
INV_X1 i_263 (.ZN (n_199), .A (n_200));
OAI21_X1 i_262 (.ZN (n_198), .A (n_201), .B1 (n_244), .B2 (n_200));
AOI21_X1 i_261 (.ZN (n_197), .A (n_198), .B1 (p_0[47]), .B2 (acc_out[47]));
NAND2_X1 i_260 (.ZN (n_196), .A1 (p_0[40]), .A2 (acc_out[40]));
NAND2_X1 i_259 (.ZN (n_195), .A1 (p_0[41]), .A2 (acc_out[41]));
INV_X1 i_258 (.ZN (n_194), .A (n_195));
AOI21_X1 i_257 (.ZN (n_193), .A (n_232), .B1 (n_196), .B2 (n_195));
AND2_X1 i_256 (.ZN (n_192), .A1 (p_0[42]), .A2 (acc_out[42]));
AOI221_X1 i_255 (.ZN (n_191), .A (n_193), .B1 (p_0[43]), .B2 (acc_out[43]), .C1 (n_237), .C2 (n_192));
OAI221_X1 i_254 (.ZN (n_190), .A (n_197), .B1 (n_239), .B2 (n_191), .C1 (n_229), .C2 (n_205));
NOR3_X1 i_253 (.ZN (n_189), .A1 (n_211), .A2 (n_190), .A3 (n_218));
NOR2_X1 i_252 (.ZN (n_188), .A1 (p_0[51]), .A2 (acc_out[51]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (p_0[49]), .A2 (acc_out[49]));
NOR2_X1 i_250 (.ZN (n_186), .A1 (p_0[50]), .A2 (acc_out[50]));
OR3_X1 i_249 (.ZN (n_185), .A1 (n_188), .A2 (n_186), .A3 (n_187));
NOR2_X1 i_248 (.ZN (n_184), .A1 (p_0[48]), .A2 (acc_out[48]));
NOR3_X1 i_247 (.ZN (n_183), .A1 (n_185), .A2 (n_184), .A3 (n_189));
NAND2_X1 i_246 (.ZN (n_182), .A1 (p_0[48]), .A2 (acc_out[48]));
NAND2_X1 i_245 (.ZN (n_181), .A1 (p_0[49]), .A2 (acc_out[49]));
AOI21_X1 i_244 (.ZN (n_180), .A (n_185), .B1 (n_182), .B2 (n_181));
AND2_X1 i_243 (.ZN (n_179), .A1 (p_0[51]), .A2 (acc_out[51]));
NAND2_X1 i_242 (.ZN (n_178), .A1 (p_0[50]), .A2 (acc_out[50]));
INV_X1 i_241 (.ZN (n_177), .A (n_178));
NOR2_X1 i_240 (.ZN (n_176), .A1 (n_188), .A2 (n_178));
NOR4_X1 i_239 (.ZN (n_175), .A1 (n_179), .A2 (n_176), .A3 (n_180), .A4 (n_183));
NOR2_X1 i_238 (.ZN (n_174), .A1 (p_0[59]), .A2 (acc_out[59]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (p_0[57]), .A2 (acc_out[57]));
NOR2_X1 i_236 (.ZN (n_172), .A1 (p_0[58]), .A2 (acc_out[58]));
NOR2_X1 i_235 (.ZN (n_171), .A1 (n_173), .A2 (n_172));
NOR3_X1 i_234 (.ZN (n_170), .A1 (n_174), .A2 (n_172), .A3 (n_173));
OAI21_X1 i_233 (.ZN (n_169), .A (n_170), .B1 (p_0[56]), .B2 (acc_out[56]));
NOR2_X1 i_232 (.ZN (n_168), .A1 (p_0[55]), .A2 (acc_out[55]));
INV_X1 i_231 (.ZN (n_167), .A (n_168));
NOR2_X1 i_230 (.ZN (n_166), .A1 (p_0[53]), .A2 (acc_out[53]));
INV_X1 i_229 (.ZN (n_165), .A (n_166));
NOR2_X1 i_228 (.ZN (n_164), .A1 (p_0[54]), .A2 (acc_out[54]));
INV_X1 i_227 (.ZN (n_163), .A (n_164));
NAND3_X1 i_226 (.ZN (n_162), .A1 (n_167), .A2 (n_163), .A3 (n_165));
NOR2_X1 i_225 (.ZN (n_161), .A1 (p_0[52]), .A2 (acc_out[52]));
OR2_X1 i_224 (.ZN (n_160), .A1 (n_162), .A2 (n_161));
NOR3_X1 i_223 (.ZN (n_159), .A1 (n_169), .A2 (n_160), .A3 (n_175));
NAND2_X1 i_222 (.ZN (n_158), .A1 (p_0[52]), .A2 (acc_out[52]));
NAND2_X1 i_221 (.ZN (n_157), .A1 (p_0[53]), .A2 (acc_out[53]));
INV_X1 i_220 (.ZN (n_156), .A (n_157));
AOI21_X1 i_219 (.ZN (n_155), .A (n_162), .B1 (n_158), .B2 (n_157));
AND2_X1 i_218 (.ZN (n_154), .A1 (p_0[54]), .A2 (acc_out[54]));
AOI221_X1 i_217 (.ZN (n_153), .A (n_155), .B1 (p_0[55]), .B2 (acc_out[55]), .C1 (n_167), .C2 (n_154));
NOR2_X1 i_216 (.ZN (n_152), .A1 (n_169), .A2 (n_153));
NAND2_X1 i_215 (.ZN (n_151), .A1 (p_0[56]), .A2 (acc_out[56]));
INV_X1 i_214 (.ZN (n_150), .A (n_151));
AND2_X1 i_213 (.ZN (n_149), .A1 (p_0[57]), .A2 (acc_out[57]));
OAI21_X1 i_212 (.ZN (n_148), .A (n_170), .B1 (n_150), .B2 (n_149));
INV_X1 i_211 (.ZN (n_147), .A (n_148));
NAND2_X1 i_210 (.ZN (n_146), .A1 (p_0[58]), .A2 (acc_out[58]));
INV_X1 i_209 (.ZN (n_145), .A (n_146));
OAI22_X1 i_208 (.ZN (n_144), .A1 (n_378), .A2 (n_374), .B1 (n_174), .B2 (n_146));
NOR4_X1 i_207 (.ZN (n_143), .A1 (n_147), .A2 (n_144), .A3 (n_152), .A4 (n_159));
AOI21_X1 i_206 (.ZN (n_142), .A (n_371), .B1 (p_0[60]), .B2 (acc_out[60]));
AOI21_X1 i_205 (.ZN (n_141), .A (n_371), .B1 (n_143), .B2 (n_142));
INV_X1 i_204 (.ZN (n_140), .A (n_141));
NAND2_X1 i_203 (.ZN (n_139), .A1 (p_0[62]), .A2 (acc_out[62]));
INV_X1 i_202 (.ZN (n_138), .A (n_139));
NAND2_X1 i_201 (.ZN (n_137), .A1 (n_379), .A2 (n_375));
OAI21_X1 i_200 (.ZN (n_136), .A (n_137), .B1 (n_379), .B2 (n_375));
INV_X1 i_199 (.ZN (n_135), .A (n_136));
NAND3_X1 i_198 (.ZN (n_134), .A1 (n_139), .A2 (n_135), .A3 (n_140));
OAI221_X1 i_197 (.ZN (n_133), .A (n_134), .B1 (p_0[62]), .B2 (acc_out[62]), .C1 (n_138), .C2 (n_137));
XNOR2_X1 i_196 (.ZN (n_132), .A (p_0[63]), .B (acc_out[63]));
XOR2_X1 i_195 (.Z (acc_out1[63]), .A (n_133), .B (n_132));
OAI21_X1 i_194 (.ZN (n_131), .A (n_139), .B1 (p_0[62]), .B2 (acc_out[62]));
AOI22_X1 i_193 (.ZN (n_130), .A1 (p_0[61]), .A2 (acc_out[61]), .B1 (n_141), .B2 (n_137));
XOR2_X1 i_192 (.Z (acc_out1[62]), .A (n_131), .B (n_130));
AOI22_X1 i_191 (.ZN (acc_out1[61]), .A1 (n_140), .A2 (n_136), .B1 (n_141), .B2 (n_135));
XNOR2_X1 i_190 (.ZN (acc_out1[60]), .A (n_143), .B (n_142));
AOI21_X1 i_189 (.ZN (n_129), .A (n_174), .B1 (p_0[59]), .B2 (acc_out[59]));
OAI21_X1 i_188 (.ZN (n_128), .A (n_153), .B1 (n_175), .B2 (n_160));
OAI21_X1 i_187 (.ZN (n_127), .A (n_151), .B1 (p_0[56]), .B2 (acc_out[56]));
OAI22_X1 i_186 (.ZN (n_126), .A1 (p_0[56]), .A2 (acc_out[56]), .B1 (n_150), .B2 (n_128));
INV_X1 i_185 (.ZN (n_125), .A (n_126));
NOR2_X1 i_184 (.ZN (n_124), .A1 (n_173), .A2 (n_149));
NAND3_X1 i_183 (.ZN (n_123), .A1 (n_146), .A2 (n_124), .A3 (n_126));
OAI21_X1 i_182 (.ZN (n_122), .A (n_123), .B1 (n_171), .B2 (n_145));
XNOR2_X1 i_181 (.ZN (acc_out1[59]), .A (n_129), .B (n_122));
NOR2_X1 i_180 (.ZN (n_121), .A1 (n_172), .A2 (n_145));
OAI22_X1 i_179 (.ZN (n_120), .A1 (p_0[57]), .A2 (acc_out[57]), .B1 (n_149), .B2 (n_125));
XNOR2_X1 i_178 (.ZN (acc_out1[58]), .A (n_121), .B (n_120));
XOR2_X1 i_177 (.Z (acc_out1[57]), .A (n_125), .B (n_124));
XNOR2_X1 i_176 (.ZN (acc_out1[56]), .A (n_128), .B (n_127));
AOI21_X1 i_175 (.ZN (n_119), .A (n_168), .B1 (p_0[55]), .B2 (acc_out[55]));
OAI21_X1 i_174 (.ZN (n_118), .A (n_158), .B1 (p_0[52]), .B2 (acc_out[52]));
AOI21_X1 i_173 (.ZN (n_117), .A (n_161), .B1 (n_175), .B2 (n_158));
OAI21_X1 i_172 (.ZN (n_116), .A (n_165), .B1 (n_156), .B2 (n_117));
INV_X1 i_171 (.ZN (n_115), .A (n_116));
NOR2_X1 i_170 (.ZN (n_114), .A1 (n_166), .A2 (n_156));
OAI21_X1 i_169 (.ZN (n_113), .A (n_163), .B1 (n_154), .B2 (n_115));
XNOR2_X1 i_168 (.ZN (acc_out1[55]), .A (n_119), .B (n_113));
NOR2_X1 i_167 (.ZN (n_112), .A1 (n_164), .A2 (n_154));
XOR2_X1 i_166 (.Z (acc_out1[54]), .A (n_115), .B (n_112));
XOR2_X1 i_165 (.Z (acc_out1[53]), .A (n_117), .B (n_114));
XOR2_X1 i_164 (.Z (acc_out1[52]), .A (n_175), .B (n_118));
NOR2_X1 i_163 (.ZN (n_111), .A1 (n_188), .A2 (n_179));
OAI21_X1 i_162 (.ZN (n_110), .A (n_182), .B1 (p_0[48]), .B2 (acc_out[48]));
AOI21_X1 i_161 (.ZN (n_109), .A (n_184), .B1 (n_189), .B2 (n_182));
INV_X1 i_160 (.ZN (n_108), .A (n_109));
AOI21_X1 i_159 (.ZN (n_107), .A (n_187), .B1 (n_181), .B2 (n_108));
AOI21_X1 i_158 (.ZN (n_106), .A (n_187), .B1 (p_0[49]), .B2 (acc_out[49]));
OAI22_X1 i_157 (.ZN (n_105), .A1 (p_0[50]), .A2 (acc_out[50]), .B1 (n_177), .B2 (n_107));
XNOR2_X1 i_156 (.ZN (acc_out1[51]), .A (n_111), .B (n_105));
NOR2_X1 i_155 (.ZN (n_104), .A1 (n_186), .A2 (n_177));
XOR2_X1 i_154 (.Z (acc_out1[50]), .A (n_107), .B (n_104));
XOR2_X1 i_153 (.Z (acc_out1[49]), .A (n_109), .B (n_106));
XOR2_X1 i_152 (.Z (acc_out1[48]), .A (n_189), .B (n_110));
AOI21_X1 i_151 (.ZN (n_103), .A (n_244), .B1 (p_0[47]), .B2 (acc_out[47]));
OAI21_X1 i_150 (.ZN (n_102), .A (n_212), .B1 (n_254), .B2 (n_219));
INV_X1 i_149 (.ZN (n_101), .A (n_102));
OAI21_X1 i_148 (.ZN (n_100), .A (n_205), .B1 (n_245), .B2 (n_101));
INV_X1 i_147 (.ZN (n_99), .A (n_100));
OAI21_X1 i_146 (.ZN (n_98), .A (n_191), .B1 (n_230), .B2 (n_99));
OAI21_X1 i_145 (.ZN (n_97), .A (n_204), .B1 (p_0[44]), .B2 (acc_out[44]));
OAI22_X1 i_144 (.ZN (n_96), .A1 (p_0[44]), .A2 (acc_out[44]), .B1 (n_203), .B2 (n_98));
INV_X1 i_143 (.ZN (n_95), .A (n_96));
NOR2_X1 i_142 (.ZN (n_94), .A1 (n_243), .A2 (n_202));
NAND3_X1 i_141 (.ZN (n_93), .A1 (n_200), .A2 (n_94), .A3 (n_96));
OAI21_X1 i_140 (.ZN (n_92), .A (n_93), .B1 (n_241), .B2 (n_199));
XNOR2_X1 i_139 (.ZN (acc_out1[47]), .A (n_103), .B (n_92));
NOR2_X1 i_138 (.ZN (n_91), .A1 (n_242), .A2 (n_199));
OAI22_X1 i_137 (.ZN (n_90), .A1 (p_0[45]), .A2 (acc_out[45]), .B1 (n_202), .B2 (n_95));
XNOR2_X1 i_136 (.ZN (acc_out1[46]), .A (n_91), .B (n_90));
XOR2_X1 i_135 (.Z (acc_out1[45]), .A (n_95), .B (n_94));
XNOR2_X1 i_134 (.ZN (acc_out1[44]), .A (n_98), .B (n_97));
AOI21_X1 i_133 (.ZN (n_89), .A (n_238), .B1 (p_0[43]), .B2 (acc_out[43]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_196), .B1 (p_0[40]), .B2 (acc_out[40]));
AOI21_X1 i_131 (.ZN (n_87), .A (n_231), .B1 (n_196), .B2 (n_99));
OAI21_X1 i_130 (.ZN (n_86), .A (n_235), .B1 (n_194), .B2 (n_87));
INV_X1 i_129 (.ZN (n_85), .A (n_86));
NOR2_X1 i_128 (.ZN (n_84), .A1 (n_236), .A2 (n_194));
OAI21_X1 i_127 (.ZN (n_83), .A (n_233), .B1 (n_192), .B2 (n_85));
XNOR2_X1 i_126 (.ZN (acc_out1[43]), .A (n_89), .B (n_83));
NOR2_X1 i_125 (.ZN (n_82), .A1 (n_234), .A2 (n_192));
XOR2_X1 i_124 (.Z (acc_out1[42]), .A (n_85), .B (n_82));
XOR2_X1 i_123 (.Z (acc_out1[41]), .A (n_87), .B (n_84));
XOR2_X1 i_122 (.Z (acc_out1[40]), .A (n_99), .B (n_88));
AOI21_X1 i_121 (.ZN (n_81), .A (n_252), .B1 (p_0[39]), .B2 (acc_out[39]));
OAI21_X1 i_120 (.ZN (n_80), .A (n_210), .B1 (p_0[36]), .B2 (acc_out[36]));
AOI21_X1 i_119 (.ZN (n_79), .A (n_253), .B1 (n_210), .B2 (n_101));
OAI21_X1 i_118 (.ZN (n_78), .A (n_249), .B1 (n_208), .B2 (n_79));
INV_X1 i_117 (.ZN (n_77), .A (n_78));
NOR2_X1 i_116 (.ZN (n_76), .A1 (n_250), .A2 (n_208));
OAI21_X1 i_115 (.ZN (n_75), .A (n_247), .B1 (n_206), .B2 (n_77));
XNOR2_X1 i_114 (.ZN (acc_out1[39]), .A (n_81), .B (n_75));
NOR2_X1 i_113 (.ZN (n_74), .A1 (n_248), .A2 (n_206));
XOR2_X1 i_112 (.Z (acc_out1[38]), .A (n_77), .B (n_74));
XOR2_X1 i_111 (.Z (acc_out1[37]), .A (n_79), .B (n_76));
XOR2_X1 i_110 (.Z (acc_out1[36]), .A (n_101), .B (n_80));
AOI21_X1 i_109 (.ZN (n_73), .A (n_227), .B1 (p_0[35]), .B2 (acc_out[35]));
OAI21_X1 i_108 (.ZN (n_72), .A (n_217), .B1 (p_0[32]), .B2 (acc_out[32]));
AOI21_X1 i_107 (.ZN (n_71), .A (n_220), .B1 (n_254), .B2 (n_217));
OAI21_X1 i_106 (.ZN (n_70), .A (n_224), .B1 (n_215), .B2 (n_71));
INV_X1 i_105 (.ZN (n_69), .A (n_70));
NOR2_X1 i_104 (.ZN (n_68), .A1 (n_225), .A2 (n_215));
OAI21_X1 i_103 (.ZN (n_67), .A (n_222), .B1 (n_213), .B2 (n_69));
XNOR2_X1 i_102 (.ZN (acc_out1[35]), .A (n_73), .B (n_67));
NOR2_X1 i_101 (.ZN (n_66), .A1 (n_223), .A2 (n_213));
XOR2_X1 i_100 (.Z (acc_out1[34]), .A (n_69), .B (n_66));
XOR2_X1 i_99 (.Z (acc_out1[33]), .A (n_71), .B (n_68));
XOR2_X1 i_98 (.Z (acc_out1[32]), .A (n_254), .B (n_72));
OAI21_X1 i_97 (.ZN (n_65), .A (n_308), .B1 (n_377), .B2 (n_373));
OAI21_X1 i_96 (.ZN (n_64), .A (n_274), .B1 (n_319), .B2 (n_281));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
OAI21_X1 i_94 (.ZN (n_62), .A (n_256), .B1 (n_310), .B2 (n_63));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
OAI21_X1 i_92 (.ZN (n_60), .A (n_268), .B1 (n_292), .B2 (n_61));
INV_X1 i_91 (.ZN (n_59), .A (n_60));
OAI21_X1 i_90 (.ZN (n_58), .A (n_267), .B1 (p_0[28]), .B2 (acc_out[28]));
AOI21_X1 i_89 (.ZN (n_57), .A (n_302), .B1 (n_267), .B2 (n_59));
OAI21_X1 i_88 (.ZN (n_56), .A (n_306), .B1 (n_266), .B2 (n_57));
INV_X1 i_87 (.ZN (n_55), .A (n_56));
NOR2_X1 i_86 (.ZN (n_54), .A1 (n_307), .A2 (n_266));
OAI21_X1 i_85 (.ZN (n_53), .A (n_304), .B1 (n_263), .B2 (n_55));
XOR2_X1 i_84 (.Z (acc_out1[31]), .A (n_65), .B (n_53));
NOR2_X1 i_83 (.ZN (n_52), .A1 (n_305), .A2 (n_263));
XOR2_X1 i_82 (.Z (acc_out1[30]), .A (n_55), .B (n_52));
XOR2_X1 i_81 (.Z (acc_out1[29]), .A (n_57), .B (n_54));
XOR2_X1 i_80 (.Z (acc_out1[28]), .A (n_59), .B (n_58));
AOI21_X1 i_79 (.ZN (n_51), .A (n_300), .B1 (p_0[27]), .B2 (acc_out[27]));
OAI21_X1 i_78 (.ZN (n_50), .A (n_273), .B1 (p_0[24]), .B2 (acc_out[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_293), .B1 (n_273), .B2 (n_61));
OAI21_X1 i_76 (.ZN (n_48), .A (n_297), .B1 (n_271), .B2 (n_49));
INV_X1 i_75 (.ZN (n_47), .A (n_48));
NOR2_X1 i_74 (.ZN (n_46), .A1 (n_298), .A2 (n_271));
OAI21_X1 i_73 (.ZN (n_45), .A (n_295), .B1 (n_269), .B2 (n_47));
XNOR2_X1 i_72 (.ZN (acc_out1[27]), .A (n_51), .B (n_45));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_296), .A2 (n_269));
XOR2_X1 i_70 (.Z (acc_out1[26]), .A (n_47), .B (n_44));
XOR2_X1 i_69 (.Z (acc_out1[25]), .A (n_49), .B (n_46));
XOR2_X1 i_68 (.Z (acc_out1[24]), .A (n_61), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_317), .B1 (p_0[23]), .B2 (acc_out[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_261), .B1 (p_0[20]), .B2 (acc_out[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_318), .B1 (n_261), .B2 (n_63));
OAI21_X1 i_64 (.ZN (n_40), .A (n_314), .B1 (n_259), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_315), .A2 (n_259));
OAI21_X1 i_61 (.ZN (n_37), .A (n_312), .B1 (n_257), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (acc_out1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_313), .A2 (n_257));
XOR2_X1 i_58 (.Z (acc_out1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (acc_out1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (acc_out1[20]), .A (n_63), .B (n_42));
AOI21_X1 i_55 (.ZN (n_35), .A (n_289), .B1 (p_0[19]), .B2 (acc_out[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_279), .B1 (p_0[16]), .B2 (acc_out[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_282), .B1 (n_319), .B2 (n_279));
OAI21_X1 i_52 (.ZN (n_32), .A (n_286), .B1 (n_277), .B2 (n_33));
INV_X1 i_51 (.ZN (n_31), .A (n_32));
NOR2_X1 i_50 (.ZN (n_30), .A1 (n_287), .A2 (n_277));
OAI21_X1 i_49 (.ZN (n_29), .A (n_284), .B1 (n_275), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (acc_out1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_285), .A2 (n_275));
XOR2_X1 i_46 (.Z (acc_out1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (acc_out1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (acc_out1[16]), .A (n_319), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_332), .A2 (n_323));
OAI21_X1 i_42 (.ZN (n_26), .A (n_326), .B1 (p_0[12]), .B2 (acc_out[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_328), .B1 (n_333), .B2 (n_326));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_331), .B1 (n_325), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_331), .B1 (p_0[13]), .B2 (acc_out[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (acc_out[14]), .B1 (n_321), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (acc_out1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_330), .A2 (n_321));
XOR2_X1 i_34 (.Z (acc_out1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (acc_out1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (acc_out1[12]), .A (n_333), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_346), .A2 (n_337));
AOI21_X1 i_30 (.ZN (n_18), .A (n_342), .B1 (p_0[8]), .B2 (acc_out[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_342), .B1 (n_347), .B2 (n_340));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_345), .B1 (n_339), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_345), .B1 (p_0[9]), .B2 (acc_out[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (acc_out[10]), .B1 (n_335), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (acc_out1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_344), .A2 (n_335));
XOR2_X1 i_22 (.Z (acc_out1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (acc_out1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (acc_out1[8]), .A (n_347), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_360), .A2 (n_351));
OAI21_X1 i_18 (.ZN (n_10), .A (n_354), .B1 (p_0[4]), .B2 (acc_out[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_356), .B1 (n_361), .B2 (n_354));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_359), .B1 (n_353), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_359), .B1 (p_0[5]), .B2 (acc_out[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (acc_out[6]), .B1 (n_349), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (acc_out1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_358), .A2 (n_349));
XOR2_X1 i_10 (.Z (acc_out1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (acc_out1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (acc_out1[4]), .A (n_361), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_370), .B1 (n_376), .B2 (n_372));
XOR2_X1 i_6 (.Z (acc_out1[3]), .A (n_363), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_369), .B1 (p_0[2]), .B2 (acc_out[2]));
XNOR2_X1 i_4 (.ZN (acc_out1[2]), .A (n_364), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_365), .B1 (p_0[1]), .B2 (acc_out[1]));
XOR2_X1 i_2 (.Z (acc_out1[1]), .A (n_366), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_366), .B1 (p_0[0]), .B2 (acc_out[0]));
INV_X1 i_0 (.ZN (acc_out1[0]), .A (n_0));

endmodule //datapath__0_10

module datapath__0_5 (p_0, in2);

output [31:0] p_0;
input [31:0] in2;
wire n_62;
wire n_60;
wire n_61;
wire n_58;
wire n_59;
wire n_5;
wire n_57;
wire n_3;
wire n_4;
wire n_1;
wire n_2;
wire n_55;
wire n_0;
wire n_56;
wire n_11;
wire n_54;
wire n_9;
wire n_10;
wire n_7;
wire n_8;
wire n_52;
wire n_6;
wire n_53;
wire n_17;
wire n_51;
wire n_15;
wire n_16;
wire n_13;
wire n_14;
wire n_49;
wire n_12;
wire n_50;
wire n_23;
wire n_48;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_45;
wire n_18;
wire n_46;
wire n_25;
wire n_44;
wire n_27;
wire n_24;
wire n_43;
wire n_26;
wire n_41;
wire n_42;
wire n_29;
wire n_40;
wire n_28;
wire n_30;
wire n_63;
wire n_32;
wire n_39;
wire n_31;
wire n_47;
wire n_34;
wire n_38;
wire n_36;
wire n_33;
wire n_37;
wire n_35;


INV_X1 i_94 (.ZN (n_63), .A (in2[25]));
NOR2_X1 i_93 (.ZN (n_62), .A1 (in2[1]), .A2 (in2[0]));
INV_X1 i_92 (.ZN (n_61), .A (n_62));
NOR2_X1 i_91 (.ZN (n_60), .A1 (in2[2]), .A2 (n_61));
INV_X1 i_90 (.ZN (n_59), .A (n_60));
NOR2_X1 i_89 (.ZN (n_58), .A1 (in2[3]), .A2 (n_59));
INV_X1 i_88 (.ZN (n_57), .A (n_58));
OR3_X1 i_87 (.ZN (n_56), .A1 (in2[6]), .A2 (in2[5]), .A3 (in2[4]));
NOR3_X1 i_86 (.ZN (n_55), .A1 (in2[7]), .A2 (n_56), .A3 (n_57));
INV_X1 i_85 (.ZN (n_54), .A (n_55));
OR3_X1 i_84 (.ZN (n_53), .A1 (in2[10]), .A2 (in2[9]), .A3 (in2[8]));
NOR3_X1 i_83 (.ZN (n_52), .A1 (in2[11]), .A2 (n_53), .A3 (n_54));
INV_X1 i_82 (.ZN (n_51), .A (n_52));
OR3_X1 i_81 (.ZN (n_50), .A1 (in2[14]), .A2 (in2[13]), .A3 (in2[12]));
NOR3_X1 i_80 (.ZN (n_49), .A1 (in2[15]), .A2 (n_50), .A3 (n_51));
INV_X1 i_79 (.ZN (n_48), .A (n_49));
OR3_X1 i_78 (.ZN (n_47), .A1 (in2[26]), .A2 (in2[25]), .A3 (in2[24]));
OR3_X1 i_77 (.ZN (n_46), .A1 (in2[18]), .A2 (in2[16]), .A3 (in2[17]));
NOR3_X1 i_76 (.ZN (n_45), .A1 (in2[19]), .A2 (n_46), .A3 (n_48));
INV_X1 i_75 (.ZN (n_44), .A (n_45));
NOR4_X1 i_74 (.ZN (n_43), .A1 (in2[22]), .A2 (in2[21]), .A3 (in2[20]), .A4 (n_44));
INV_X1 i_73 (.ZN (n_42), .A (n_43));
NOR2_X1 i_72 (.ZN (n_41), .A1 (in2[23]), .A2 (n_42));
INV_X1 i_71 (.ZN (n_40), .A (n_41));
NOR3_X1 i_70 (.ZN (n_39), .A1 (in2[27]), .A2 (n_47), .A3 (n_40));
INV_X1 i_69 (.ZN (n_38), .A (n_39));
NOR4_X1 i_68 (.ZN (n_37), .A1 (in2[29]), .A2 (in2[28]), .A3 (in2[30]), .A4 (n_38));
XNOR2_X1 i_67 (.ZN (p_0[31]), .A (in2[31]), .B (n_37));
NOR3_X1 i_66 (.ZN (n_36), .A1 (in2[29]), .A2 (in2[28]), .A3 (n_38));
INV_X1 i_65 (.ZN (n_35), .A (n_36));
AOI21_X1 i_64 (.ZN (p_0[30]), .A (n_37), .B1 (in2[30]), .B2 (n_35));
NOR2_X1 i_63 (.ZN (n_34), .A1 (in2[28]), .A2 (n_38));
INV_X1 i_62 (.ZN (n_33), .A (n_34));
AOI21_X1 i_61 (.ZN (p_0[29]), .A (n_36), .B1 (in2[29]), .B2 (n_33));
AOI21_X1 i_60 (.ZN (p_0[28]), .A (n_34), .B1 (in2[28]), .B2 (n_38));
NOR2_X1 i_59 (.ZN (n_32), .A1 (n_47), .A2 (n_40));
INV_X1 i_58 (.ZN (n_31), .A (n_32));
AOI21_X1 i_57 (.ZN (p_0[27]), .A (n_39), .B1 (in2[27]), .B2 (n_31));
OR3_X1 i_56 (.ZN (n_30), .A1 (in2[25]), .A2 (in2[24]), .A3 (n_40));
AOI21_X1 i_55 (.ZN (p_0[26]), .A (n_32), .B1 (in2[26]), .B2 (n_30));
NOR2_X1 i_54 (.ZN (n_29), .A1 (in2[24]), .A2 (n_40));
OAI21_X1 i_53 (.ZN (n_28), .A (n_30), .B1 (n_63), .B2 (n_29));
INV_X1 i_52 (.ZN (p_0[25]), .A (n_28));
AOI21_X1 i_51 (.ZN (p_0[24]), .A (n_29), .B1 (in2[24]), .B2 (n_40));
AOI21_X1 i_50 (.ZN (p_0[23]), .A (n_41), .B1 (in2[23]), .B2 (n_42));
NOR3_X1 i_49 (.ZN (n_27), .A1 (in2[21]), .A2 (in2[20]), .A3 (n_44));
INV_X1 i_48 (.ZN (n_26), .A (n_27));
AOI21_X1 i_47 (.ZN (p_0[22]), .A (n_43), .B1 (in2[22]), .B2 (n_26));
NOR2_X1 i_46 (.ZN (n_25), .A1 (in2[20]), .A2 (n_44));
INV_X1 i_45 (.ZN (n_24), .A (n_25));
AOI21_X1 i_44 (.ZN (p_0[21]), .A (n_27), .B1 (in2[21]), .B2 (n_24));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_25), .B1 (in2[20]), .B2 (n_44));
NOR2_X1 i_42 (.ZN (n_23), .A1 (in2[16]), .A2 (n_48));
INV_X1 i_41 (.ZN (n_22), .A (n_23));
NOR2_X1 i_40 (.ZN (n_21), .A1 (in2[17]), .A2 (n_22));
INV_X1 i_39 (.ZN (n_20), .A (n_21));
NOR2_X1 i_38 (.ZN (n_19), .A1 (n_48), .A2 (n_46));
INV_X1 i_37 (.ZN (n_18), .A (n_19));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_45), .B1 (in2[19]), .B2 (n_18));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_19), .B1 (in2[18]), .B2 (n_20));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_21), .B1 (in2[17]), .B2 (n_22));
AOI21_X1 i_33 (.ZN (p_0[16]), .A (n_23), .B1 (in2[16]), .B2 (n_48));
NOR2_X1 i_32 (.ZN (n_17), .A1 (in2[12]), .A2 (n_51));
INV_X1 i_31 (.ZN (n_16), .A (n_17));
NOR2_X1 i_30 (.ZN (n_15), .A1 (in2[13]), .A2 (n_16));
INV_X1 i_29 (.ZN (n_14), .A (n_15));
NOR2_X1 i_28 (.ZN (n_13), .A1 (n_51), .A2 (n_50));
INV_X1 i_27 (.ZN (n_12), .A (n_13));
AOI21_X1 i_26 (.ZN (p_0[15]), .A (n_49), .B1 (in2[15]), .B2 (n_12));
AOI21_X1 i_25 (.ZN (p_0[14]), .A (n_13), .B1 (in2[14]), .B2 (n_14));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_15), .B1 (in2[13]), .B2 (n_16));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_17), .B1 (in2[12]), .B2 (n_51));
NOR2_X1 i_22 (.ZN (n_11), .A1 (in2[8]), .A2 (n_54));
INV_X1 i_21 (.ZN (n_10), .A (n_11));
NOR2_X1 i_20 (.ZN (n_9), .A1 (in2[9]), .A2 (n_10));
INV_X1 i_19 (.ZN (n_8), .A (n_9));
NOR2_X1 i_18 (.ZN (n_7), .A1 (n_54), .A2 (n_53));
INV_X1 i_17 (.ZN (n_6), .A (n_7));
AOI21_X1 i_16 (.ZN (p_0[11]), .A (n_52), .B1 (in2[11]), .B2 (n_6));
AOI21_X1 i_15 (.ZN (p_0[10]), .A (n_7), .B1 (in2[10]), .B2 (n_8));
AOI21_X1 i_14 (.ZN (p_0[9]), .A (n_9), .B1 (in2[9]), .B2 (n_10));
AOI21_X1 i_13 (.ZN (p_0[8]), .A (n_11), .B1 (in2[8]), .B2 (n_54));
NOR2_X1 i_12 (.ZN (n_5), .A1 (in2[4]), .A2 (n_57));
INV_X1 i_11 (.ZN (n_4), .A (n_5));
NOR2_X1 i_10 (.ZN (n_3), .A1 (in2[5]), .A2 (n_4));
INV_X1 i_9 (.ZN (n_2), .A (n_3));
NOR2_X1 i_8 (.ZN (n_1), .A1 (n_57), .A2 (n_56));
INV_X1 i_7 (.ZN (n_0), .A (n_1));
AOI21_X1 i_6 (.ZN (p_0[7]), .A (n_55), .B1 (in2[7]), .B2 (n_0));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_1), .B1 (in2[6]), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_0[5]), .A (n_3), .B1 (in2[5]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (in2[4]), .B2 (n_57));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_58), .B1 (in2[3]), .B2 (n_59));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_60), .B1 (in2[2]), .B2 (n_61));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_62), .B1 (in2[1]), .B2 (in2[0]));

endmodule //datapath__0_5

module datapath (p_0, in1);

output [31:0] p_0;
input [31:0] in1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (in1[25]));
INV_X1 i_63 (.ZN (n_32), .A (in1[21]));
INV_X1 i_62 (.ZN (n_31), .A (in1[14]));
INV_X1 i_61 (.ZN (n_30), .A (in1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (in1[2]), .A2 (in1[1]), .A3 (in1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (in1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (in1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (in1[5]), .A3 (in1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (in1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (in1[8]), .A3 (in1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (in1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (in1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (in1[12]), .A3 (in1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (in1[15]), .A3 (in1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (in1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (in1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (in1[18]), .A3 (in1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (in1[18]), .A3 (in1[19]), .A4 (in1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (in1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (in1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (in1[23]), .A3 (in1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (in1[26]), .A3 (in1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (in1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (in1[28]), .A3 (in1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (in1[28]), .A3 (in1[29]), .A4 (in1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (in1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (in1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (in1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (in1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (in1[27]), .B1 (n_9), .B2 (in1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (in1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (in1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (in1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (in1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (in1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (in1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (in1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (in1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (in1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (in1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (in1[16]), .B1 (n_19), .B2 (in1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (in1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (in1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (in1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (in1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (in1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (in1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (in1[9]), .B1 (n_25), .B2 (in1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (in1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (in1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (in1[6]), .B1 (n_27), .B2 (in1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (in1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (in1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (in1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (in1[2]), .B1 (in1[1]), .B2 (in1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (in1[1]), .B (in1[0]));

endmodule //datapath

module sequential_multiplier (clk_CTSPP_233, clk_CTSPP_229, clk_CTSPP_230, clk_CTSPP_231, 
    clk_CTSPP_234, clk_CTSPP_236, clk, rst, in1, in2, out);

output [63:0] out;
output clk_CTSPP_233;
input clk;
input [31:0] in1;
input [31:0] in2;
input rst;
input clk_CTSPP_229;
input clk_CTSPP_230;
input clk_CTSPP_231;
input clk_CTSPP_234;
input clk_CTSPP_236;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire n_0_317;
wire n_0_318;
wire n_0_319;
wire n_0_320;
wire n_0_321;
wire n_0_322;
wire n_0_323;
wire n_0_324;
wire n_0_325;
wire n_0_326;
wire n_0_327;
wire n_0_328;
wire n_0_329;
wire n_0_330;
wire n_0_331;
wire n_0_332;
wire n_0_333;
wire n_0_334;
wire n_0_335;
wire n_0_336;
wire n_0_337;
wire n_0_338;
wire n_0_339;
wire n_0_340;
wire n_0_341;
wire n_0_342;
wire n_0_343;
wire n_0_344;
wire n_0_345;
wire n_0_346;
wire n_0_347;
wire n_0_348;
wire n_0_349;
wire n_0_350;
wire n_0_351;
wire n_0_352;
wire n_0_353;
wire n_0_354;
wire n_0_355;
wire n_0_356;
wire n_0_357;
wire n_0_358;
wire n_0_359;
wire n_0_360;
wire n_0_361;
wire n_0_362;
wire n_0_363;
wire n_0_364;
wire n_0_365;
wire n_0_366;
wire n_0_367;
wire n_0_368;
wire n_0_369;
wire n_0_370;
wire n_0_371;
wire n_0_372;
wire n_0_373;
wire n_0_374;
wire n_0_375;
wire n_0_376;
wire n_0_377;
wire n_0_378;
wire n_0_379;
wire n_0_380;
wire n_0_381;
wire n_0_382;
wire n_0_383;
wire n_0_384;
wire n_0_385;
wire n_0_386;
wire n_0_387;
wire n_0_388;
wire n_0_389;
wire n_0_390;
wire n_0_391;
wire n_0_392;
wire n_0_393;
wire n_0_394;
wire n_0_395;
wire n_0_396;
wire n_0_397;
wire n_0_398;
wire n_0_399;
wire n_0_400;
wire n_0_401;
wire n_0_402;
wire n_0_403;
wire n_0_404;
wire n_0_405;
wire n_0_406;
wire n_0_407;
wire n_0_408;
wire n_0_409;
wire n_0_410;
wire n_0_411;
wire n_0_412;
wire n_0_413;
wire n_0_414;
wire n_0_415;
wire n_0_416;
wire n_0_417;
wire n_0_418;
wire n_0_419;
wire n_0_420;
wire n_0_421;
wire n_0_422;
wire n_0_423;
wire n_0_424;
wire n_0_425;
wire n_0_426;
wire n_0_427;
wire n_0_428;
wire n_0_429;
wire n_0_430;
wire n_0_431;
wire n_0_432;
wire n_0_433;
wire n_0_434;
wire n_0_435;
wire n_0_436;
wire n_0_437;
wire n_0_438;
wire n_0_439;
wire n_0_440;
wire n_0_441;
wire n_0_442;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire \A1[63] ;
wire \A1[62] ;
wire \A1[61] ;
wire \A1[60] ;
wire \A1[59] ;
wire \A1[58] ;
wire \A1[57] ;
wire \A1[56] ;
wire \A1[55] ;
wire \A1[54] ;
wire \A1[53] ;
wire \A1[52] ;
wire \A1[51] ;
wire \A1[50] ;
wire \A1[49] ;
wire \A1[48] ;
wire \A1[47] ;
wire \A1[46] ;
wire \A1[45] ;
wire \A1[44] ;
wire \A1[43] ;
wire \A1[42] ;
wire \A1[41] ;
wire \A1[40] ;
wire \A1[39] ;
wire \A1[38] ;
wire \A1[37] ;
wire \A1[36] ;
wire \A1[35] ;
wire \A1[34] ;
wire \A1[33] ;
wire \A1[32] ;
wire \A1[31] ;
wire \A1[30] ;
wire \A1[29] ;
wire \A1[28] ;
wire \A1[27] ;
wire \A1[26] ;
wire \A1[25] ;
wire \A1[24] ;
wire \A1[23] ;
wire \A1[22] ;
wire \A1[21] ;
wire \A1[20] ;
wire \A1[19] ;
wire \A1[18] ;
wire \A1[17] ;
wire \A1[16] ;
wire \A1[15] ;
wire \A1[14] ;
wire \A1[13] ;
wire \A1[12] ;
wire \A1[11] ;
wire \A1[10] ;
wire \A1[9] ;
wire \A1[8] ;
wire \A1[7] ;
wire \A1[6] ;
wire \A1[5] ;
wire \A1[4] ;
wire \A1[3] ;
wire \A1[2] ;
wire \A1[1] ;
wire \A1[0] ;
wire \B1[31] ;
wire \B1[30] ;
wire \B1[29] ;
wire \B1[28] ;
wire \B1[27] ;
wire \B1[26] ;
wire \B1[25] ;
wire \B1[24] ;
wire \B1[23] ;
wire \B1[22] ;
wire \B1[21] ;
wire \B1[20] ;
wire \B1[19] ;
wire \B1[18] ;
wire \B1[17] ;
wire \B1[16] ;
wire \B1[15] ;
wire \B1[14] ;
wire \B1[13] ;
wire \B1[12] ;
wire \B1[11] ;
wire \B1[10] ;
wire \B1[9] ;
wire \B1[8] ;
wire \B1[7] ;
wire \B1[6] ;
wire \B1[5] ;
wire \B1[4] ;
wire \B1[3] ;
wire \B1[2] ;
wire \B1[1] ;
wire \B1[0] ;
wire \acc_out[63] ;
wire \acc_out[62] ;
wire \acc_out[61] ;
wire \acc_out[60] ;
wire \acc_out[59] ;
wire \acc_out[58] ;
wire \acc_out[57] ;
wire \acc_out[56] ;
wire \acc_out[55] ;
wire \acc_out[54] ;
wire \acc_out[53] ;
wire \acc_out[52] ;
wire \acc_out[51] ;
wire \acc_out[50] ;
wire \acc_out[49] ;
wire \acc_out[48] ;
wire \acc_out[47] ;
wire \acc_out[46] ;
wire \acc_out[45] ;
wire \acc_out[44] ;
wire \acc_out[43] ;
wire \acc_out[42] ;
wire \acc_out[41] ;
wire \acc_out[40] ;
wire \acc_out[39] ;
wire \acc_out[38] ;
wire \acc_out[37] ;
wire \acc_out[36] ;
wire \acc_out[35] ;
wire \acc_out[34] ;
wire \acc_out[33] ;
wire \acc_out[32] ;
wire \acc_out[31] ;
wire \acc_out[30] ;
wire \acc_out[29] ;
wire \acc_out[28] ;
wire \acc_out[27] ;
wire \acc_out[26] ;
wire \acc_out[25] ;
wire \acc_out[24] ;
wire \acc_out[23] ;
wire \acc_out[22] ;
wire \acc_out[21] ;
wire \acc_out[20] ;
wire \acc_out[19] ;
wire \acc_out[18] ;
wire \acc_out[17] ;
wire \acc_out[16] ;
wire \acc_out[15] ;
wire \acc_out[14] ;
wire \acc_out[13] ;
wire \acc_out[12] ;
wire \acc_out[11] ;
wire \acc_out[10] ;
wire \acc_out[9] ;
wire \acc_out[8] ;
wire \acc_out[7] ;
wire \acc_out[6] ;
wire \acc_out[5] ;
wire \acc_out[4] ;
wire \acc_out[3] ;
wire \acc_out[2] ;
wire \acc_out[1] ;
wire \acc_out[0] ;
wire n_354;
wire CTS_n105;
wire n_193;
wire n_192;
wire n_191;
wire n_190;
wire n_189;
wire n_188;
wire n_187;
wire n_186;
wire n_185;
wire n_184;
wire n_183;
wire n_182;
wire n_181;
wire n_180;
wire n_179;
wire n_178;
wire n_177;
wire n_176;
wire n_175;
wire n_174;
wire n_173;
wire n_172;
wire n_171;
wire n_170;
wire n_169;
wire n_168;
wire n_167;
wire n_166;
wire n_165;
wire n_164;
wire n_163;
wire n_162;
wire n_161;
wire n_160;
wire n_159;
wire n_158;
wire n_157;
wire n_156;
wire n_155;
wire n_154;
wire n_153;
wire n_152;
wire n_151;
wire n_150;
wire n_149;
wire n_148;
wire n_147;
wire n_146;
wire n_145;
wire n_144;
wire n_143;
wire n_142;
wire n_141;
wire n_140;
wire n_139;
wire n_138;
wire n_137;
wire n_136;
wire n_135;
wire n_134;
wire n_133;
wire n_132;
wire n_131;
wire n_130;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire uc_0;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire uc_1;
wire n_321;
wire n_320;
wire n_319;
wire n_318;
wire n_317;
wire n_316;
wire n_315;
wire n_314;
wire n_313;
wire n_312;
wire n_311;
wire n_310;
wire n_309;
wire n_308;
wire n_307;
wire n_306;
wire n_305;
wire n_304;
wire n_303;
wire n_302;
wire n_301;
wire n_300;
wire n_299;
wire n_298;
wire n_297;
wire n_296;
wire n_295;
wire n_294;
wire n_293;
wire n_292;
wire n_291;
wire n_290;
wire n_289;
wire n_288;
wire n_287;
wire n_286;
wire n_285;
wire n_284;
wire n_283;
wire n_282;
wire n_281;
wire n_280;
wire n_279;
wire n_278;
wire n_277;
wire n_276;
wire n_275;
wire n_274;
wire n_273;
wire n_272;
wire n_271;
wire n_270;
wire n_269;
wire n_268;
wire n_267;
wire n_266;
wire n_265;
wire n_264;
wire n_263;
wire n_262;
wire n_261;
wire n_260;
wire n_259;
wire n_258;
wire n_257;
wire n_256;
wire n_255;
wire n_254;
wire n_253;
wire n_252;
wire n_251;
wire n_250;
wire n_249;
wire n_248;
wire n_247;
wire n_246;
wire n_245;
wire n_244;
wire n_243;
wire n_242;
wire n_241;
wire n_240;
wire n_239;
wire n_238;
wire n_237;
wire n_236;
wire n_235;
wire n_234;
wire n_233;
wire n_232;
wire n_231;
wire n_230;
wire n_229;
wire n_228;
wire n_227;
wire n_226;
wire n_225;
wire n_224;
wire n_223;
wire n_222;
wire n_221;
wire n_220;
wire n_219;
wire n_218;
wire n_217;
wire n_216;
wire n_215;
wire n_214;
wire n_213;
wire n_212;
wire n_211;
wire n_210;
wire n_209;
wire n_208;
wire n_207;
wire n_206;
wire n_205;
wire n_204;
wire n_203;
wire n_202;
wire n_201;
wire n_200;
wire n_199;
wire n_198;
wire n_197;
wire n_196;
wire n_195;
wire n_194;
wire n_126;
wire n_125;
wire n_124;
wire n_123;
wire n_122;
wire n_121;
wire n_120;
wire n_119;
wire n_118;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_104;
wire n_103;
wire n_102;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_127;
wire n_128;
wire n_129;
wire n_355;
wire n_357;
wire n_327;
wire n_326;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_356;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire hfn_ipo_n72;
wire hfn_ipo_n73;
wire hfn_ipo_n71;
wire hfn_ipo_n74;
wire hfn_ipo_n76;
wire hfn_ipo_n77;
wire hfn_ipo_n75;
wire hfn_ipo_n78;
wire hfn_ipo_n79;
wire hfn_ipo_n80;
wire hfn_ipo_n82;
wire hfn_ipo_n83;
wire hfn_ipo_n81;
wire CTS_n106;
wire hfn_ipo_n94;
wire hfn_ipo_n95;
wire hfn_ipo_n86;
wire hfn_ipo_n87;
wire hfn_ipo_n85;
wire hfn_ipo_n88;
wire hfn_ipo_n89;
wire hfn_ipo_n90;
wire hfn_ipo_n91;
wire hfn_ipo_n92;
wire hfn_ipo_n65;
wire hfn_ipo_n66;
wire hfn_ipo_n67;
wire hfn_ipo_n68;
wire hfn_ipo_n69;
wire drc_ipo_n96;
wire hfn_ipo_n70;
wire CLOCK_slh__n1277;


DFF_X1 \acc_out_reg[0]  (.Q (\acc_out[0] ), .CK (clk_CTSPP_233), .D (n_63));
DFF_X1 \acc_out_reg[1]  (.Q (\acc_out[1] ), .CK (clk_CTSPP_233), .D (n_64));
DFF_X1 \acc_out_reg[2]  (.Q (\acc_out[2] ), .CK (clk_CTSPP_233), .D (n_65));
DFF_X1 \acc_out_reg[3]  (.Q (\acc_out[3] ), .CK (clk_CTSPP_233), .D (n_66));
DFF_X1 \acc_out_reg[4]  (.Q (\acc_out[4] ), .CK (clk_CTSPP_233), .D (n_67));
DFF_X1 \acc_out_reg[5]  (.Q (\acc_out[5] ), .CK (clk_CTSPP_233), .D (n_68));
DFF_X1 \acc_out_reg[6]  (.Q (\acc_out[6] ), .CK (clk_CTSPP_234), .D (n_69));
DFF_X1 \acc_out_reg[7]  (.Q (\acc_out[7] ), .CK (clk_CTSPP_234), .D (n_70));
DFF_X1 \acc_out_reg[8]  (.Q (\acc_out[8] ), .CK (clk_CTSPP_234), .D (n_71));
DFF_X1 \acc_out_reg[9]  (.Q (\acc_out[9] ), .CK (clk_CTSPP_234), .D (n_72));
DFF_X1 \acc_out_reg[10]  (.Q (\acc_out[10] ), .CK (clk_CTSPP_234), .D (n_73));
DFF_X1 \acc_out_reg[11]  (.Q (\acc_out[11] ), .CK (clk_CTSPP_234), .D (n_74));
DFF_X1 \acc_out_reg[12]  (.Q (\acc_out[12] ), .CK (clk_CTSPP_234), .D (n_75));
DFF_X1 \acc_out_reg[13]  (.Q (\acc_out[13] ), .CK (clk_CTSPP_234), .D (n_76));
DFF_X1 \acc_out_reg[14]  (.Q (\acc_out[14] ), .CK (clk_CTSPP_234), .D (n_77));
DFF_X1 \acc_out_reg[15]  (.Q (\acc_out[15] ), .CK (clk_CTSPP_234), .D (n_78));
DFF_X1 \acc_out_reg[16]  (.Q (\acc_out[16] ), .CK (clk_CTSPP_233), .D (n_79));
DFF_X1 \acc_out_reg[17]  (.Q (\acc_out[17] ), .CK (clk_CTSPP_234), .D (n_80));
DFF_X1 \acc_out_reg[18]  (.Q (\acc_out[18] ), .CK (clk_CTSPP_234), .D (n_81));
DFF_X1 \acc_out_reg[19]  (.Q (\acc_out[19] ), .CK (clk_CTSPP_234), .D (n_82));
DFF_X1 \acc_out_reg[20]  (.Q (\acc_out[20] ), .CK (clk_CTSPP_234), .D (n_83));
DFF_X1 \acc_out_reg[21]  (.Q (\acc_out[21] ), .CK (clk_CTSPP_233), .D (n_84));
DFF_X1 \acc_out_reg[22]  (.Q (\acc_out[22] ), .CK (clk_CTSPP_233), .D (n_85));
DFF_X1 \acc_out_reg[23]  (.Q (\acc_out[23] ), .CK (clk_CTSPP_233), .D (n_86));
DFF_X1 \acc_out_reg[24]  (.Q (\acc_out[24] ), .CK (clk_CTSPP_233), .D (n_87));
DFF_X1 \acc_out_reg[25]  (.Q (\acc_out[25] ), .CK (clk_CTSPP_233), .D (n_88));
DFF_X1 \acc_out_reg[26]  (.Q (\acc_out[26] ), .CK (clk_CTSPP_233), .D (n_89));
DFF_X1 \acc_out_reg[27]  (.Q (\acc_out[27] ), .CK (clk_CTSPP_233), .D (n_90));
DFF_X1 \acc_out_reg[28]  (.Q (\acc_out[28] ), .CK (clk_CTSPP_233), .D (n_91));
DFF_X1 \acc_out_reg[29]  (.Q (\acc_out[29] ), .CK (clk_CTSPP_233), .D (n_92));
DFF_X1 \acc_out_reg[30]  (.Q (\acc_out[30] ), .CK (clk_CTSPP_233), .D (n_93));
DFF_X1 \acc_out_reg[31]  (.Q (\acc_out[31] ), .CK (clk_CTSPP_234), .D (n_94));
DFF_X1 \acc_out_reg[32]  (.Q (\acc_out[32] ), .CK (clk_CTSPP_234), .D (n_95));
DFF_X1 \acc_out_reg[33]  (.Q (\acc_out[33] ), .CK (clk_CTSPP_233), .D (n_96));
DFF_X1 \acc_out_reg[34]  (.Q (\acc_out[34] ), .CK (clk_CTSPP_234), .D (n_97));
DFF_X1 \acc_out_reg[35]  (.Q (\acc_out[35] ), .CK (clk_CTSPP_234), .D (n_98));
DFF_X1 \acc_out_reg[36]  (.Q (\acc_out[36] ), .CK (clk_CTSPP_234), .D (n_99));
DFF_X1 \acc_out_reg[37]  (.Q (\acc_out[37] ), .CK (clk_CTSPP_234), .D (n_100));
DFF_X1 \acc_out_reg[38]  (.Q (\acc_out[38] ), .CK (clk_CTSPP_234), .D (n_101));
DFF_X1 \acc_out_reg[39]  (.Q (\acc_out[39] ), .CK (clk_CTSPP_234), .D (n_102));
DFF_X1 \acc_out_reg[40]  (.Q (\acc_out[40] ), .CK (clk_CTSPP_234), .D (n_103));
DFF_X1 \acc_out_reg[41]  (.Q (\acc_out[41] ), .CK (clk_CTSPP_234), .D (n_104));
DFF_X1 \acc_out_reg[42]  (.Q (\acc_out[42] ), .CK (clk_CTSPP_234), .D (n_105));
DFF_X1 \acc_out_reg[43]  (.Q (\acc_out[43] ), .CK (clk_CTSPP_234), .D (n_106));
DFF_X1 \acc_out_reg[44]  (.Q (\acc_out[44] ), .CK (clk_CTSPP_234), .D (n_107));
DFF_X1 \acc_out_reg[45]  (.Q (\acc_out[45] ), .CK (clk_CTSPP_230), .D (n_108));
DFF_X1 \acc_out_reg[46]  (.Q (\acc_out[46] ), .CK (clk_CTSPP_230), .D (n_109));
DFF_X1 \acc_out_reg[47]  (.Q (\acc_out[47] ), .CK (clk_CTSPP_234), .D (n_110));
DFF_X1 \acc_out_reg[48]  (.Q (\acc_out[48] ), .CK (clk_CTSPP_230), .D (n_111));
DFF_X1 \acc_out_reg[49]  (.Q (\acc_out[49] ), .CK (clk_CTSPP_230), .D (n_112));
DFF_X1 \acc_out_reg[50]  (.Q (\acc_out[50] ), .CK (clk_CTSPP_230), .D (n_113));
DFF_X1 \acc_out_reg[51]  (.Q (\acc_out[51] ), .CK (clk_CTSPP_230), .D (n_114));
DFF_X1 \acc_out_reg[52]  (.Q (\acc_out[52] ), .CK (clk_CTSPP_230), .D (n_115));
DFF_X1 \acc_out_reg[53]  (.Q (\acc_out[53] ), .CK (clk_CTSPP_230), .D (n_116));
DFF_X1 \acc_out_reg[54]  (.Q (\acc_out[54] ), .CK (clk_CTSPP_230), .D (n_117));
DFF_X1 \acc_out_reg[55]  (.Q (\acc_out[55] ), .CK (clk_CTSPP_230), .D (n_118));
DFF_X1 \acc_out_reg[56]  (.Q (\acc_out[56] ), .CK (clk_CTSPP_230), .D (n_119));
DFF_X1 \acc_out_reg[57]  (.Q (\acc_out[57] ), .CK (clk_CTSPP_230), .D (n_120));
DFF_X1 \acc_out_reg[58]  (.Q (\acc_out[58] ), .CK (clk_CTSPP_230), .D (n_121));
DFF_X1 \acc_out_reg[59]  (.Q (\acc_out[59] ), .CK (clk_CTSPP_230), .D (n_122));
DFF_X1 \acc_out_reg[60]  (.Q (\acc_out[60] ), .CK (clk_CTSPP_230), .D (n_123));
DFF_X1 \acc_out_reg[61]  (.Q (\acc_out[61] ), .CK (clk_CTSPP_230), .D (n_124));
DFF_X1 \acc_out_reg[62]  (.Q (\acc_out[62] ), .CK (clk_CTSPP_230), .D (n_125));
DFF_X1 \acc_out_reg[63]  (.Q (\acc_out[63] ), .CK (clk_CTSPP_230), .D (n_126));
DFF_X1 \B1_reg[0]  (.Q (\B1[0] ), .CK (clk_CTSPP_229), .D (n_322));
DFF_X1 \B1_reg[1]  (.Q (\B1[1] ), .CK (clk_CTSPP_229), .D (n_323));
DFF_X1 \B1_reg[2]  (.Q (\B1[2] ), .CK (clk_CTSPP_229), .D (n_324));
DFF_X1 \B1_reg[3]  (.Q (\B1[3] ), .CK (clk_CTSPP_229), .D (n_325));
DFF_X1 \B1_reg[4]  (.Q (\B1[4] ), .CK (clk_CTSPP_229), .D (n_326));
DFF_X1 \B1_reg[5]  (.Q (\B1[5] ), .CK (clk_CTSPP_229), .D (n_327));
DFF_X1 \B1_reg[6]  (.Q (\B1[6] ), .CK (clk_CTSPP_229), .D (n_328));
DFF_X1 \B1_reg[7]  (.Q (\B1[7] ), .CK (clk_CTSPP_229), .D (n_329));
DFF_X1 \B1_reg[8]  (.Q (\B1[8] ), .CK (clk_CTSPP_229), .D (n_330));
DFF_X1 \B1_reg[9]  (.Q (\B1[9] ), .CK (clk_CTSPP_233), .D (n_331));
DFF_X1 \B1_reg[10]  (.Q (\B1[10] ), .CK (clk_CTSPP_229), .D (n_332));
DFF_X1 \B1_reg[11]  (.Q (\B1[11] ), .CK (clk_CTSPP_229), .D (n_333));
DFF_X1 \B1_reg[12]  (.Q (\B1[12] ), .CK (clk_CTSPP_229), .D (n_334));
DFF_X1 \B1_reg[13]  (.Q (\B1[13] ), .CK (clk_CTSPP_233), .D (n_335));
DFF_X1 \B1_reg[14]  (.Q (\B1[14] ), .CK (clk_CTSPP_229), .D (n_336));
DFF_X1 \B1_reg[15]  (.Q (\B1[15] ), .CK (clk_CTSPP_229), .D (n_337));
DFF_X1 \B1_reg[16]  (.Q (\B1[16] ), .CK (clk_CTSPP_229), .D (n_338));
DFF_X1 \B1_reg[17]  (.Q (\B1[17] ), .CK (clk_CTSPP_229), .D (n_339));
DFF_X1 \B1_reg[18]  (.Q (\B1[18] ), .CK (clk_CTSPP_229), .D (n_340));
DFF_X1 \B1_reg[19]  (.Q (\B1[19] ), .CK (clk_CTSPP_229), .D (n_341));
DFF_X1 \B1_reg[20]  (.Q (\B1[20] ), .CK (clk_CTSPP_229), .D (n_342));
DFF_X1 \B1_reg[21]  (.Q (\B1[21] ), .CK (clk_CTSPP_229), .D (n_343));
DFF_X1 \B1_reg[22]  (.Q (\B1[22] ), .CK (clk_CTSPP_229), .D (n_344));
DFF_X1 \B1_reg[23]  (.Q (\B1[23] ), .CK (clk_CTSPP_229), .D (n_345));
DFF_X1 \B1_reg[24]  (.Q (\B1[24] ), .CK (clk_CTSPP_231), .D (n_346));
DFF_X1 \B1_reg[25]  (.Q (\B1[25] ), .CK (clk_CTSPP_229), .D (n_347));
DFF_X1 \B1_reg[26]  (.Q (\B1[26] ), .CK (clk_CTSPP_229), .D (n_348));
DFF_X1 \B1_reg[27]  (.Q (\B1[27] ), .CK (clk_CTSPP_229), .D (n_349));
DFF_X1 \B1_reg[28]  (.Q (\B1[28] ), .CK (clk_CTSPP_231), .D (n_350));
DFF_X1 \B1_reg[29]  (.Q (\B1[29] ), .CK (clk_CTSPP_231), .D (n_351));
DFF_X1 \B1_reg[30]  (.Q (\B1[30] ), .CK (clk_CTSPP_229), .D (n_352));
DFF_X1 \B1_reg[31]  (.Q (\B1[31] ), .CK (clk_CTSPP_229), .D (n_353));
DFF_X1 \A1_reg[0]  (.Q (\A1[0] ), .CK (clk_CTSPP_233), .D (n_357));
DFF_X1 \A1_reg[1]  (.Q (\A1[1] ), .CK (clk_CTSPP_233), .D (n_358));
DFF_X1 \A1_reg[2]  (.Q (\A1[2] ), .CK (clk_CTSPP_233), .D (n_359));
DFF_X1 \A1_reg[3]  (.Q (\A1[3] ), .CK (clk_CTSPP_229), .D (n_360));
DFF_X1 \A1_reg[4]  (.Q (\A1[4] ), .CK (clk_CTSPP_229), .D (n_361));
DFF_X1 \A1_reg[5]  (.Q (\A1[5] ), .CK (clk_CTSPP_229), .D (n_362));
DFF_X1 \A1_reg[6]  (.Q (\A1[6] ), .CK (clk_CTSPP_229), .D (n_363));
DFF_X1 \A1_reg[7]  (.Q (\A1[7] ), .CK (clk_CTSPP_233), .D (n_364));
DFF_X1 \A1_reg[8]  (.Q (\A1[8] ), .CK (clk_CTSPP_233), .D (n_365));
DFF_X1 \A1_reg[9]  (.Q (\A1[9] ), .CK (clk_CTSPP_233), .D (n_366));
DFF_X1 \A1_reg[10]  (.Q (\A1[10] ), .CK (clk_CTSPP_231), .D (n_367));
DFF_X1 \A1_reg[11]  (.Q (\A1[11] ), .CK (clk_CTSPP_231), .D (n_368));
DFF_X1 \A1_reg[12]  (.Q (\A1[12] ), .CK (clk_CTSPP_231), .D (n_369));
DFF_X1 \A1_reg[13]  (.Q (\A1[13] ), .CK (clk_CTSPP_231), .D (n_370));
DFF_X1 \A1_reg[14]  (.Q (\A1[14] ), .CK (clk_CTSPP_231), .D (n_371));
DFF_X1 \A1_reg[15]  (.Q (\A1[15] ), .CK (clk_CTSPP_231), .D (n_372));
DFF_X1 \A1_reg[16]  (.Q (\A1[16] ), .CK (clk_CTSPP_231), .D (n_373));
DFF_X1 \A1_reg[17]  (.Q (\A1[17] ), .CK (clk_CTSPP_229), .D (n_374));
DFF_X1 \A1_reg[18]  (.Q (\A1[18] ), .CK (clk_CTSPP_229), .D (n_375));
DFF_X1 \A1_reg[19]  (.Q (\A1[19] ), .CK (clk_CTSPP_229), .D (n_376));
DFF_X1 \A1_reg[20]  (.Q (\A1[20] ), .CK (clk_CTSPP_229), .D (n_377));
DFF_X1 \A1_reg[21]  (.Q (\A1[21] ), .CK (clk_CTSPP_231), .D (n_378));
DFF_X1 \A1_reg[22]  (.Q (\A1[22] ), .CK (clk_CTSPP_231), .D (n_379));
DFF_X1 \A1_reg[23]  (.Q (\A1[23] ), .CK (clk_CTSPP_231), .D (n_380));
DFF_X1 \A1_reg[24]  (.Q (\A1[24] ), .CK (clk_CTSPP_231), .D (n_381));
DFF_X1 \A1_reg[25]  (.Q (\A1[25] ), .CK (clk_CTSPP_231), .D (n_382));
DFF_X1 \A1_reg[26]  (.Q (\A1[26] ), .CK (clk_CTSPP_230), .D (n_383));
DFF_X1 \A1_reg[27]  (.Q (\A1[27] ), .CK (clk_CTSPP_231), .D (n_384));
DFF_X1 \A1_reg[28]  (.Q (\A1[28] ), .CK (clk_CTSPP_230), .D (n_385));
DFF_X1 \A1_reg[29]  (.Q (\A1[29] ), .CK (clk_CTSPP_230), .D (n_386));
DFF_X1 \A1_reg[30]  (.Q (\A1[30] ), .CK (clk_CTSPP_230), .D (n_387));
DFF_X1 \A1_reg[31]  (.Q (\A1[31] ), .CK (clk_CTSPP_231), .D (n_388));
DFF_X1 \A1_reg[32]  (.Q (\A1[32] ), .CK (clk_CTSPP_231), .D (n_389));
DFF_X1 \A1_reg[33]  (.Q (\A1[33] ), .CK (clk_CTSPP_231), .D (n_390));
DFF_X1 \A1_reg[34]  (.Q (\A1[34] ), .CK (clk_CTSPP_231), .D (n_391));
DFF_X1 \A1_reg[35]  (.Q (\A1[35] ), .CK (clk_CTSPP_231), .D (n_392));
DFF_X1 \A1_reg[36]  (.Q (\A1[36] ), .CK (clk_CTSPP_231), .D (n_393));
DFF_X1 \A1_reg[37]  (.Q (\A1[37] ), .CK (clk_CTSPP_230), .D (n_394));
DFF_X1 \A1_reg[38]  (.Q (\A1[38] ), .CK (clk_CTSPP_230), .D (n_395));
DFF_X1 \A1_reg[39]  (.Q (\A1[39] ), .CK (clk_CTSPP_231), .D (n_396));
DFF_X1 \A1_reg[40]  (.Q (\A1[40] ), .CK (clk_CTSPP_231), .D (n_397));
DFF_X1 \A1_reg[41]  (.Q (\A1[41] ), .CK (clk_CTSPP_231), .D (n_398));
DFF_X1 \A1_reg[42]  (.Q (\A1[42] ), .CK (clk_CTSPP_230), .D (n_399));
DFF_X1 \A1_reg[43]  (.Q (\A1[43] ), .CK (clk_CTSPP_230), .D (n_400));
DFF_X1 \A1_reg[44]  (.Q (\A1[44] ), .CK (clk_CTSPP_231), .D (n_401));
DFF_X1 \A1_reg[45]  (.Q (\A1[45] ), .CK (clk_CTSPP_231), .D (n_402));
DFF_X1 \A1_reg[46]  (.Q (\A1[46] ), .CK (clk_CTSPP_231), .D (n_403));
DFF_X1 \A1_reg[47]  (.Q (\A1[47] ), .CK (clk_CTSPP_231), .D (n_404));
DFF_X1 \A1_reg[48]  (.Q (\A1[48] ), .CK (clk_CTSPP_231), .D (n_405));
DFF_X1 \A1_reg[49]  (.Q (\A1[49] ), .CK (clk_CTSPP_231), .D (n_406));
DFF_X1 \A1_reg[50]  (.Q (\A1[50] ), .CK (clk_CTSPP_230), .D (n_407));
DFF_X1 \A1_reg[51]  (.Q (\A1[51] ), .CK (clk_CTSPP_231), .D (n_408));
DFF_X1 \A1_reg[52]  (.Q (\A1[52] ), .CK (clk_CTSPP_231), .D (n_409));
DFF_X1 \A1_reg[53]  (.Q (\A1[53] ), .CK (clk_CTSPP_230), .D (n_410));
DFF_X1 \A1_reg[54]  (.Q (\A1[54] ), .CK (clk_CTSPP_230), .D (n_411));
DFF_X1 \A1_reg[55]  (.Q (\A1[55] ), .CK (clk_CTSPP_231), .D (n_412));
DFF_X1 \A1_reg[56]  (.Q (\A1[56] ), .CK (clk_CTSPP_231), .D (n_413));
DFF_X1 \A1_reg[57]  (.Q (\A1[57] ), .CK (clk_CTSPP_230), .D (n_414));
DFF_X1 \A1_reg[58]  (.Q (\A1[58] ), .CK (clk_CTSPP_230), .D (n_415));
DFF_X1 \A1_reg[59]  (.Q (\A1[59] ), .CK (clk_CTSPP_230), .D (n_416));
DFF_X1 \A1_reg[60]  (.Q (\A1[60] ), .CK (clk_CTSPP_231), .D (n_417));
DFF_X1 \A1_reg[61]  (.Q (\A1[61] ), .CK (clk_CTSPP_230), .D (n_418));
DFF_X1 \A1_reg[62]  (.Q (\A1[62] ), .CK (clk_CTSPP_230), .D (n_419));
DFF_X1 \A1_reg[63]  (.Q (\A1[63] ), .CK (clk_CTSPP_230), .D (n_420));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (clk_CTSPP_229), .D (hfn_ipo_n94));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (clk_CTSPP_229), .D (n_127));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (clk_CTSPP_229), .D (n_128));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (clk_CTSPP_229), .D (n_129));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (clk_CTSPP_229), .D (n_356));
INV_X1 i_0_733 (.ZN (n_0_442), .A (rst));
INV_X1 i_0_732 (.ZN (n_0_441), .A (in1[31]));
INV_X1 i_0_731 (.ZN (n_0_440), .A (\counter[0] ));
INV_X1 i_0_730 (.ZN (n_0_439), .A (\A1[0] ));
NOR2_X1 i_0_729 (.ZN (n_0_438), .A1 (hfn_ipo_n89), .A2 (in2[31]));
AND2_X1 i_0_728 (.ZN (n_0_437), .A1 (in1[31]), .A2 (hfn_ipo_n88));
AND2_X1 i_0_727 (.ZN (n_0_436), .A1 (rst), .A2 (in2[31]));
AOI221_X1 i_0_726 (.ZN (n_0_435), .A (n_0_437), .B1 (n_0_441), .B2 (hfn_ipo_n86), .C1 (n_31), .C2 (hfn_ipo_n86));
INV_X2 i_0_725 (.ZN (n_0_434), .A (n_0_435));
AOI21_X1 i_0_724 (.ZN (n_0_433), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[63] ));
INV_X1 i_0_723 (.ZN (n_420), .A (n_0_433));
AOI21_X1 i_0_722 (.ZN (n_0_432), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[62] ));
INV_X1 i_0_721 (.ZN (n_419), .A (n_0_432));
AOI21_X1 i_0_720 (.ZN (n_0_431), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[61] ));
INV_X1 i_0_719 (.ZN (n_418), .A (n_0_431));
AOI21_X1 i_0_718 (.ZN (n_0_430), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[60] ));
INV_X1 i_0_717 (.ZN (n_417), .A (n_0_430));
AOI21_X1 i_0_716 (.ZN (n_0_429), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[59] ));
INV_X1 i_0_715 (.ZN (n_416), .A (n_0_429));
AOI21_X1 i_0_714 (.ZN (n_0_428), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[58] ));
INV_X1 i_0_713 (.ZN (n_415), .A (n_0_428));
AOI21_X1 i_0_712 (.ZN (n_0_427), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[57] ));
INV_X1 i_0_711 (.ZN (n_414), .A (n_0_427));
AOI21_X1 i_0_710 (.ZN (n_0_426), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[56] ));
INV_X1 i_0_709 (.ZN (n_413), .A (n_0_426));
AOI21_X1 i_0_708 (.ZN (n_0_425), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[55] ));
INV_X1 i_0_707 (.ZN (n_412), .A (n_0_425));
AOI21_X1 i_0_706 (.ZN (n_0_424), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[54] ));
INV_X1 i_0_705 (.ZN (n_411), .A (n_0_424));
AOI21_X1 i_0_704 (.ZN (n_0_423), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[53] ));
INV_X1 i_0_703 (.ZN (n_410), .A (n_0_423));
AOI21_X1 i_0_702 (.ZN (n_0_422), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[52] ));
INV_X1 i_0_701 (.ZN (n_409), .A (n_0_422));
AOI21_X1 i_0_700 (.ZN (n_0_421), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[51] ));
INV_X1 i_0_699 (.ZN (n_408), .A (n_0_421));
AOI21_X1 i_0_698 (.ZN (n_0_420), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[50] ));
INV_X1 i_0_697 (.ZN (n_407), .A (n_0_420));
AOI21_X1 i_0_696 (.ZN (n_0_419), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[49] ));
INV_X1 i_0_695 (.ZN (n_406), .A (n_0_419));
AOI21_X1 i_0_694 (.ZN (n_0_418), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[48] ));
INV_X1 i_0_693 (.ZN (n_405), .A (n_0_418));
AOI21_X1 i_0_692 (.ZN (n_0_417), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[47] ));
INV_X1 i_0_691 (.ZN (n_404), .A (n_0_417));
AOI21_X1 i_0_690 (.ZN (n_0_416), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[46] ));
INV_X1 i_0_689 (.ZN (n_403), .A (n_0_416));
AOI21_X1 i_0_688 (.ZN (n_0_415), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[45] ));
INV_X1 i_0_687 (.ZN (n_402), .A (n_0_415));
AOI21_X1 i_0_686 (.ZN (n_0_414), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[44] ));
INV_X1 i_0_685 (.ZN (n_401), .A (n_0_414));
AOI21_X1 i_0_684 (.ZN (n_0_413), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[43] ));
INV_X1 i_0_683 (.ZN (n_400), .A (n_0_413));
AOI21_X1 i_0_682 (.ZN (n_0_412), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[42] ));
INV_X1 i_0_681 (.ZN (n_399), .A (n_0_412));
AOI21_X1 i_0_680 (.ZN (n_0_411), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[41] ));
INV_X1 i_0_679 (.ZN (n_398), .A (n_0_411));
AOI21_X1 i_0_678 (.ZN (n_0_410), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[40] ));
INV_X1 i_0_677 (.ZN (n_397), .A (n_0_410));
AOI21_X1 i_0_676 (.ZN (n_0_409), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[39] ));
INV_X1 i_0_675 (.ZN (n_396), .A (n_0_409));
AOI21_X1 i_0_674 (.ZN (n_0_408), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[38] ));
INV_X1 i_0_673 (.ZN (n_395), .A (n_0_408));
AOI21_X1 i_0_672 (.ZN (n_0_407), .A (n_0_434), .B1 (n_0_442), .B2 (\A1[37] ));
INV_X1 i_0_671 (.ZN (n_394), .A (n_0_407));
AOI21_X1 i_0_670 (.ZN (n_0_406), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[36] ));
INV_X1 i_0_669 (.ZN (n_393), .A (n_0_406));
AOI21_X1 i_0_668 (.ZN (n_0_405), .A (n_0_434), .B1 (hfn_ipo_n92), .B2 (\A1[35] ));
INV_X1 i_0_667 (.ZN (n_392), .A (n_0_405));
AOI21_X1 i_0_666 (.ZN (n_0_404), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[34] ));
INV_X1 i_0_665 (.ZN (n_391), .A (n_0_404));
AOI21_X1 i_0_664 (.ZN (n_0_403), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[33] ));
INV_X1 i_0_663 (.ZN (n_390), .A (n_0_403));
AOI21_X1 i_0_662 (.ZN (n_0_402), .A (n_0_434), .B1 (hfn_ipo_n91), .B2 (\A1[32] ));
INV_X1 i_0_661 (.ZN (n_389), .A (n_0_402));
AOI221_X1 i_0_660 (.ZN (n_0_401), .A (n_0_437), .B1 (hfn_ipo_n92), .B2 (\A1[31] )
    , .C1 (n_31), .C2 (hfn_ipo_n86));
INV_X1 i_0_659 (.ZN (n_388), .A (n_0_401));
AOI222_X1 i_0_658 (.ZN (n_0_400), .A1 (hfn_ipo_n92), .A2 (\A1[30] ), .B1 (in1[30])
    , .B2 (hfn_ipo_n88), .C1 (n_30), .C2 (hfn_ipo_n86));
INV_X1 i_0_657 (.ZN (n_387), .A (n_0_400));
AOI222_X1 i_0_656 (.ZN (n_0_399), .A1 (hfn_ipo_n92), .A2 (\A1[29] ), .B1 (in1[29])
    , .B2 (hfn_ipo_n88), .C1 (n_29), .C2 (hfn_ipo_n86));
INV_X1 i_0_655 (.ZN (n_386), .A (n_0_399));
AOI222_X1 i_0_654 (.ZN (n_0_398), .A1 (hfn_ipo_n92), .A2 (\A1[28] ), .B1 (in1[28])
    , .B2 (hfn_ipo_n88), .C1 (n_28), .C2 (hfn_ipo_n86));
INV_X1 i_0_653 (.ZN (n_385), .A (n_0_398));
AOI222_X1 i_0_652 (.ZN (n_0_397), .A1 (hfn_ipo_n92), .A2 (\A1[27] ), .B1 (in1[27])
    , .B2 (hfn_ipo_n88), .C1 (n_27), .C2 (hfn_ipo_n86));
INV_X1 i_0_651 (.ZN (n_384), .A (n_0_397));
AOI222_X1 i_0_650 (.ZN (n_0_396), .A1 (hfn_ipo_n92), .A2 (\A1[26] ), .B1 (in1[26])
    , .B2 (hfn_ipo_n88), .C1 (n_26), .C2 (hfn_ipo_n86));
INV_X1 i_0_649 (.ZN (n_383), .A (n_0_396));
AOI222_X1 i_0_648 (.ZN (n_0_395), .A1 (hfn_ipo_n92), .A2 (\A1[25] ), .B1 (in1[25])
    , .B2 (hfn_ipo_n88), .C1 (n_25), .C2 (hfn_ipo_n86));
INV_X1 i_0_647 (.ZN (n_382), .A (n_0_395));
AOI222_X1 i_0_646 (.ZN (n_0_394), .A1 (hfn_ipo_n92), .A2 (\A1[24] ), .B1 (in1[24])
    , .B2 (hfn_ipo_n88), .C1 (n_24), .C2 (hfn_ipo_n86));
INV_X1 i_0_645 (.ZN (n_381), .A (n_0_394));
AOI222_X1 i_0_644 (.ZN (n_0_393), .A1 (hfn_ipo_n92), .A2 (\A1[23] ), .B1 (in1[23])
    , .B2 (hfn_ipo_n88), .C1 (n_23), .C2 (hfn_ipo_n86));
INV_X1 i_0_643 (.ZN (n_380), .A (n_0_393));
AOI222_X1 i_0_642 (.ZN (n_0_392), .A1 (hfn_ipo_n89), .A2 (\A1[22] ), .B1 (in1[22])
    , .B2 (hfn_ipo_n88), .C1 (n_22), .C2 (hfn_ipo_n86));
INV_X1 i_0_641 (.ZN (n_379), .A (n_0_392));
AOI222_X1 i_0_640 (.ZN (n_0_391), .A1 (hfn_ipo_n89), .A2 (\A1[21] ), .B1 (in1[21])
    , .B2 (hfn_ipo_n88), .C1 (n_21), .C2 (hfn_ipo_n86));
INV_X1 i_0_639 (.ZN (n_378), .A (n_0_391));
AOI222_X1 i_0_638 (.ZN (n_0_390), .A1 (hfn_ipo_n89), .A2 (\A1[20] ), .B1 (in1[20])
    , .B2 (hfn_ipo_n88), .C1 (n_20), .C2 (hfn_ipo_n86));
INV_X1 i_0_637 (.ZN (n_377), .A (n_0_390));
AOI222_X1 i_0_636 (.ZN (n_0_389), .A1 (hfn_ipo_n89), .A2 (\A1[19] ), .B1 (in1[19])
    , .B2 (hfn_ipo_n88), .C1 (n_19), .C2 (hfn_ipo_n86));
INV_X1 i_0_635 (.ZN (n_376), .A (n_0_389));
AOI222_X1 i_0_634 (.ZN (n_0_388), .A1 (hfn_ipo_n89), .A2 (\A1[18] ), .B1 (in1[18])
    , .B2 (hfn_ipo_n88), .C1 (n_18), .C2 (hfn_ipo_n86));
INV_X1 i_0_633 (.ZN (n_375), .A (n_0_388));
AOI222_X1 i_0_632 (.ZN (n_0_387), .A1 (hfn_ipo_n89), .A2 (\A1[17] ), .B1 (in1[17])
    , .B2 (hfn_ipo_n88), .C1 (n_17), .C2 (hfn_ipo_n86));
INV_X1 i_0_631 (.ZN (n_374), .A (n_0_387));
AOI222_X1 i_0_630 (.ZN (n_0_386), .A1 (hfn_ipo_n92), .A2 (\A1[16] ), .B1 (in1[16])
    , .B2 (hfn_ipo_n88), .C1 (n_16), .C2 (hfn_ipo_n86));
INV_X1 i_0_629 (.ZN (n_373), .A (n_0_386));
AOI222_X1 i_0_628 (.ZN (n_0_385), .A1 (hfn_ipo_n92), .A2 (\A1[15] ), .B1 (in1[15])
    , .B2 (hfn_ipo_n88), .C1 (n_15), .C2 (hfn_ipo_n86));
INV_X1 i_0_627 (.ZN (n_372), .A (n_0_385));
AOI222_X1 i_0_626 (.ZN (n_0_384), .A1 (hfn_ipo_n92), .A2 (\A1[14] ), .B1 (in1[14])
    , .B2 (hfn_ipo_n88), .C1 (n_14), .C2 (hfn_ipo_n86));
INV_X1 i_0_625 (.ZN (n_371), .A (n_0_384));
AOI222_X1 i_0_624 (.ZN (n_0_383), .A1 (hfn_ipo_n92), .A2 (\A1[13] ), .B1 (in1[13])
    , .B2 (hfn_ipo_n88), .C1 (n_13), .C2 (hfn_ipo_n86));
INV_X1 i_0_623 (.ZN (n_370), .A (n_0_383));
AOI222_X1 i_0_622 (.ZN (n_0_382), .A1 (hfn_ipo_n92), .A2 (\A1[12] ), .B1 (in1[12])
    , .B2 (hfn_ipo_n88), .C1 (n_12), .C2 (hfn_ipo_n86));
INV_X1 i_0_621 (.ZN (n_369), .A (n_0_382));
AOI222_X1 i_0_620 (.ZN (n_0_381), .A1 (hfn_ipo_n91), .A2 (\A1[11] ), .B1 (in1[11])
    , .B2 (hfn_ipo_n88), .C1 (n_11), .C2 (hfn_ipo_n86));
INV_X1 i_0_619 (.ZN (n_368), .A (n_0_381));
AOI222_X1 i_0_618 (.ZN (n_0_380), .A1 (hfn_ipo_n90), .A2 (\A1[10] ), .B1 (in1[10])
    , .B2 (hfn_ipo_n88), .C1 (n_10), .C2 (hfn_ipo_n86));
INV_X1 i_0_617 (.ZN (n_367), .A (n_0_380));
AOI222_X1 i_0_616 (.ZN (n_0_379), .A1 (hfn_ipo_n90), .A2 (\A1[9] ), .B1 (in1[9]), .B2 (hfn_ipo_n88)
    , .C1 (n_9), .C2 (hfn_ipo_n86));
INV_X1 i_0_615 (.ZN (n_366), .A (n_0_379));
AOI222_X1 i_0_614 (.ZN (n_0_378), .A1 (hfn_ipo_n90), .A2 (\A1[8] ), .B1 (in1[8]), .B2 (hfn_ipo_n88)
    , .C1 (n_8), .C2 (hfn_ipo_n86));
INV_X1 i_0_613 (.ZN (n_365), .A (n_0_378));
AOI222_X1 i_0_612 (.ZN (n_0_377), .A1 (hfn_ipo_n90), .A2 (\A1[7] ), .B1 (in1[7]), .B2 (hfn_ipo_n88)
    , .C1 (n_7), .C2 (hfn_ipo_n86));
INV_X1 i_0_611 (.ZN (n_364), .A (n_0_377));
AOI222_X1 i_0_610 (.ZN (n_0_376), .A1 (hfn_ipo_n90), .A2 (\A1[6] ), .B1 (in1[6]), .B2 (hfn_ipo_n87)
    , .C1 (n_6), .C2 (hfn_ipo_n85));
INV_X1 i_0_609 (.ZN (n_363), .A (n_0_376));
AOI222_X1 i_0_608 (.ZN (n_0_375), .A1 (hfn_ipo_n89), .A2 (\A1[5] ), .B1 (in1[5]), .B2 (hfn_ipo_n87)
    , .C1 (n_5), .C2 (hfn_ipo_n85));
INV_X1 i_0_607 (.ZN (n_362), .A (n_0_375));
AOI222_X1 i_0_606 (.ZN (n_0_374), .A1 (hfn_ipo_n89), .A2 (\A1[4] ), .B1 (in1[4]), .B2 (hfn_ipo_n87)
    , .C1 (n_4), .C2 (hfn_ipo_n85));
INV_X1 i_0_605 (.ZN (n_361), .A (n_0_374));
AOI222_X1 i_0_604 (.ZN (n_0_373), .A1 (hfn_ipo_n89), .A2 (\A1[3] ), .B1 (in1[3]), .B2 (hfn_ipo_n87)
    , .C1 (n_3), .C2 (hfn_ipo_n85));
INV_X1 i_0_603 (.ZN (n_360), .A (n_0_373));
AOI222_X1 i_0_602 (.ZN (n_0_372), .A1 (hfn_ipo_n90), .A2 (\A1[2] ), .B1 (in1[2]), .B2 (hfn_ipo_n87)
    , .C1 (n_2), .C2 (hfn_ipo_n85));
INV_X1 i_0_601 (.ZN (n_359), .A (n_0_372));
AOI222_X1 i_0_600 (.ZN (n_0_371), .A1 (hfn_ipo_n90), .A2 (\A1[1] ), .B1 (in1[1]), .B2 (hfn_ipo_n87)
    , .C1 (n_1), .C2 (hfn_ipo_n85));
INV_X1 i_0_599 (.ZN (n_358), .A (n_0_371));
NAND2_X1 i_0_598 (.ZN (n_0_370), .A1 (rst), .A2 (in1[0]));
OAI21_X1 i_0_597 (.ZN (n_357), .A (n_0_370), .B1 (rst), .B2 (n_0_439));
NAND2_X1 i_0_596 (.ZN (n_0_369), .A1 (hfn_ipo_n89), .A2 (\counter[4] ));
INV_X1 i_0_595 (.ZN (n_0_368), .A (hfn_ipo_n83));
XNOR2_X1 i_0_594 (.ZN (n_356), .A (n_0_2), .B (hfn_ipo_n83));
NAND2_X1 i_0_593 (.ZN (n_355), .A1 (hfn_ipo_n89), .A2 (\counter[0] ));
INV_X1 i_0_592 (.ZN (n_0_367), .A (hfn_ipo_n94));
NAND2_X1 i_0_591 (.ZN (n_0_366), .A1 (hfn_ipo_n89), .A2 (\counter[3] ));
INV_X1 i_0_590 (.ZN (n_0_365), .A (hfn_ipo_n77));
NAND4_X1 i_0_589 (.ZN (n_0_364), .A1 (\counter[1] ), .A2 (n_0_440), .A3 (\counter[4] ), .A4 (\counter[2] ));
NOR2_X1 i_0_588 (.ZN (n_0_363), .A1 (hfn_ipo_n77), .A2 (n_0_364));
OAI21_X1 i_0_587 (.ZN (n_354), .A (hfn_ipo_n89), .B1 (hfn_ipo_n77), .B2 (n_0_364));
AOI22_X1 i_0_586 (.ZN (n_0_362), .A1 (n_62), .A2 (hfn_ipo_n86), .B1 (hfn_ipo_n89), .B2 (\B1[31] ));
INV_X1 i_0_585 (.ZN (n_353), .A (n_0_362));
AOI222_X1 i_0_584 (.ZN (n_0_361), .A1 (hfn_ipo_n89), .A2 (\B1[30] ), .B1 (in2[30])
    , .B2 (hfn_ipo_n88), .C1 (n_61), .C2 (hfn_ipo_n86));
INV_X1 i_0_583 (.ZN (n_352), .A (n_0_361));
AOI222_X1 i_0_582 (.ZN (n_0_360), .A1 (hfn_ipo_n89), .A2 (\B1[29] ), .B1 (in2[29])
    , .B2 (hfn_ipo_n88), .C1 (n_60), .C2 (hfn_ipo_n86));
INV_X1 i_0_581 (.ZN (n_351), .A (n_0_360));
AOI222_X1 i_0_580 (.ZN (n_0_359), .A1 (hfn_ipo_n89), .A2 (\B1[28] ), .B1 (in2[28])
    , .B2 (hfn_ipo_n88), .C1 (n_59), .C2 (hfn_ipo_n86));
INV_X1 i_0_579 (.ZN (n_350), .A (n_0_359));
AOI222_X1 i_0_578 (.ZN (n_0_358), .A1 (hfn_ipo_n89), .A2 (\B1[27] ), .B1 (in2[27])
    , .B2 (hfn_ipo_n87), .C1 (n_58), .C2 (hfn_ipo_n85));
INV_X1 i_0_577 (.ZN (n_349), .A (n_0_358));
AOI222_X1 i_0_576 (.ZN (n_0_357), .A1 (hfn_ipo_n89), .A2 (\B1[26] ), .B1 (in2[26])
    , .B2 (hfn_ipo_n87), .C1 (n_57), .C2 (hfn_ipo_n85));
INV_X1 i_0_575 (.ZN (n_348), .A (n_0_357));
AOI222_X1 i_0_574 (.ZN (n_0_356), .A1 (hfn_ipo_n89), .A2 (\B1[25] ), .B1 (in2[25])
    , .B2 (hfn_ipo_n88), .C1 (n_56), .C2 (hfn_ipo_n85));
INV_X1 i_0_573 (.ZN (n_347), .A (n_0_356));
AOI222_X1 i_0_572 (.ZN (n_0_355), .A1 (hfn_ipo_n89), .A2 (\B1[24] ), .B1 (in2[24])
    , .B2 (hfn_ipo_n88), .C1 (n_55), .C2 (hfn_ipo_n86));
INV_X1 i_0_571 (.ZN (n_346), .A (n_0_355));
AOI222_X1 i_0_570 (.ZN (n_0_354), .A1 (hfn_ipo_n89), .A2 (\B1[23] ), .B1 (in2[23])
    , .B2 (hfn_ipo_n87), .C1 (n_54), .C2 (hfn_ipo_n85));
INV_X1 i_0_569 (.ZN (n_345), .A (n_0_354));
AOI222_X1 i_0_568 (.ZN (n_0_353), .A1 (hfn_ipo_n89), .A2 (\B1[22] ), .B1 (in2[22])
    , .B2 (hfn_ipo_n87), .C1 (n_53), .C2 (hfn_ipo_n85));
INV_X1 i_0_567 (.ZN (n_344), .A (n_0_353));
AOI222_X1 i_0_566 (.ZN (n_0_352), .A1 (hfn_ipo_n89), .A2 (\B1[21] ), .B1 (in2[21])
    , .B2 (hfn_ipo_n87), .C1 (n_52), .C2 (hfn_ipo_n85));
INV_X1 i_0_565 (.ZN (n_343), .A (n_0_352));
AOI222_X1 i_0_564 (.ZN (n_0_351), .A1 (hfn_ipo_n89), .A2 (\B1[20] ), .B1 (in2[20])
    , .B2 (hfn_ipo_n87), .C1 (n_51), .C2 (hfn_ipo_n85));
INV_X1 i_0_563 (.ZN (n_342), .A (n_0_351));
AOI222_X1 i_0_562 (.ZN (n_0_350), .A1 (hfn_ipo_n89), .A2 (\B1[19] ), .B1 (in2[19])
    , .B2 (hfn_ipo_n87), .C1 (n_50), .C2 (hfn_ipo_n85));
INV_X1 i_0_561 (.ZN (n_341), .A (n_0_350));
AOI222_X1 i_0_560 (.ZN (n_0_349), .A1 (hfn_ipo_n89), .A2 (\B1[18] ), .B1 (in2[18])
    , .B2 (hfn_ipo_n87), .C1 (n_49), .C2 (hfn_ipo_n85));
INV_X1 i_0_559 (.ZN (n_340), .A (n_0_349));
AOI222_X1 i_0_558 (.ZN (n_0_348), .A1 (hfn_ipo_n89), .A2 (\B1[17] ), .B1 (in2[17])
    , .B2 (hfn_ipo_n87), .C1 (n_48), .C2 (hfn_ipo_n85));
INV_X1 i_0_557 (.ZN (n_339), .A (n_0_348));
AOI222_X1 i_0_556 (.ZN (n_0_347), .A1 (hfn_ipo_n89), .A2 (\B1[16] ), .B1 (in2[16])
    , .B2 (hfn_ipo_n87), .C1 (n_47), .C2 (hfn_ipo_n85));
INV_X1 i_0_555 (.ZN (n_338), .A (n_0_347));
AOI222_X1 i_0_554 (.ZN (n_0_346), .A1 (hfn_ipo_n89), .A2 (\B1[15] ), .B1 (in2[15])
    , .B2 (hfn_ipo_n87), .C1 (n_46), .C2 (hfn_ipo_n85));
INV_X1 i_0_553 (.ZN (n_337), .A (n_0_346));
AOI222_X1 i_0_552 (.ZN (n_0_345), .A1 (hfn_ipo_n89), .A2 (\B1[14] ), .B1 (in2[14])
    , .B2 (hfn_ipo_n87), .C1 (n_45), .C2 (hfn_ipo_n85));
INV_X1 i_0_551 (.ZN (n_336), .A (n_0_345));
AOI222_X1 i_0_550 (.ZN (n_0_344), .A1 (hfn_ipo_n89), .A2 (\B1[13] ), .B1 (in2[13])
    , .B2 (hfn_ipo_n87), .C1 (n_44), .C2 (hfn_ipo_n85));
INV_X1 i_0_549 (.ZN (n_335), .A (n_0_344));
AOI222_X1 i_0_548 (.ZN (n_0_343), .A1 (hfn_ipo_n89), .A2 (\B1[12] ), .B1 (in2[12])
    , .B2 (hfn_ipo_n87), .C1 (n_43), .C2 (hfn_ipo_n85));
INV_X1 i_0_547 (.ZN (n_334), .A (n_0_343));
AOI222_X1 i_0_546 (.ZN (n_0_342), .A1 (hfn_ipo_n89), .A2 (\B1[11] ), .B1 (in2[11])
    , .B2 (hfn_ipo_n87), .C1 (n_42), .C2 (hfn_ipo_n85));
INV_X1 i_0_545 (.ZN (n_333), .A (n_0_342));
AOI222_X1 i_0_544 (.ZN (n_0_341), .A1 (hfn_ipo_n89), .A2 (\B1[10] ), .B1 (in2[10])
    , .B2 (hfn_ipo_n87), .C1 (n_41), .C2 (hfn_ipo_n85));
INV_X1 i_0_543 (.ZN (n_332), .A (n_0_341));
AOI222_X1 i_0_542 (.ZN (n_0_340), .A1 (hfn_ipo_n89), .A2 (\B1[9] ), .B1 (in2[9]), .B2 (hfn_ipo_n87)
    , .C1 (n_40), .C2 (hfn_ipo_n85));
INV_X1 i_0_541 (.ZN (n_331), .A (n_0_340));
AOI222_X1 i_0_540 (.ZN (n_0_339), .A1 (hfn_ipo_n89), .A2 (\B1[8] ), .B1 (in2[8]), .B2 (hfn_ipo_n87)
    , .C1 (n_39), .C2 (hfn_ipo_n85));
INV_X1 i_0_539 (.ZN (n_330), .A (n_0_339));
AOI222_X1 i_0_538 (.ZN (n_0_338), .A1 (hfn_ipo_n89), .A2 (\B1[7] ), .B1 (in2[7]), .B2 (hfn_ipo_n87)
    , .C1 (n_38), .C2 (hfn_ipo_n85));
INV_X1 i_0_537 (.ZN (n_329), .A (n_0_338));
AOI222_X1 i_0_536 (.ZN (n_0_337), .A1 (hfn_ipo_n89), .A2 (\B1[6] ), .B1 (in2[6]), .B2 (hfn_ipo_n87)
    , .C1 (n_37), .C2 (hfn_ipo_n85));
INV_X1 i_0_535 (.ZN (n_328), .A (n_0_337));
AOI222_X1 i_0_534 (.ZN (n_0_336), .A1 (hfn_ipo_n89), .A2 (\B1[5] ), .B1 (in2[5]), .B2 (hfn_ipo_n87)
    , .C1 (n_36), .C2 (hfn_ipo_n85));
INV_X1 i_0_533 (.ZN (n_327), .A (n_0_336));
AOI222_X1 i_0_532 (.ZN (n_0_335), .A1 (hfn_ipo_n89), .A2 (\B1[4] ), .B1 (in2[4]), .B2 (hfn_ipo_n87)
    , .C1 (n_35), .C2 (hfn_ipo_n85));
INV_X1 i_0_531 (.ZN (n_326), .A (n_0_335));
AOI222_X1 i_0_530 (.ZN (n_0_334), .A1 (hfn_ipo_n89), .A2 (\B1[3] ), .B1 (in2[3]), .B2 (hfn_ipo_n87)
    , .C1 (n_34), .C2 (hfn_ipo_n85));
INV_X1 i_0_529 (.ZN (n_325), .A (n_0_334));
AOI222_X1 i_0_528 (.ZN (n_0_333), .A1 (hfn_ipo_n89), .A2 (\B1[2] ), .B1 (in2[2]), .B2 (hfn_ipo_n87)
    , .C1 (n_33), .C2 (hfn_ipo_n85));
INV_X1 i_0_527 (.ZN (n_324), .A (n_0_333));
AOI222_X1 i_0_526 (.ZN (n_0_332), .A1 (hfn_ipo_n89), .A2 (\B1[1] ), .B1 (in2[1]), .B2 (hfn_ipo_n87)
    , .C1 (n_32), .C2 (hfn_ipo_n85));
INV_X1 i_0_525 (.ZN (n_323), .A (n_0_332));
AOI22_X1 i_0_524 (.ZN (n_0_331), .A1 (hfn_ipo_n89), .A2 (\B1[0] ), .B1 (rst), .B2 (in2[0]));
INV_X1 i_0_523 (.ZN (CLOCK_slh__n1277), .A (n_0_331));
NAND2_X1 i_0_522 (.ZN (n_0_330), .A1 (hfn_ipo_n89), .A2 (\counter[1] ));
INV_X1 i_0_521 (.ZN (n_0_329), .A (hfn_ipo_n72));
NAND2_X1 i_0_520 (.ZN (n_0_328), .A1 (hfn_ipo_n89), .A2 (\counter[2] ));
INV_X1 i_0_519 (.ZN (n_0_327), .A (hfn_ipo_n67));
AOI22_X1 i_0_518 (.ZN (n_0_326), .A1 (\counter[0] ), .A2 (n_0_354), .B1 (n_0_440), .B2 (n_0_353));
AOI22_X1 i_0_517 (.ZN (n_0_325), .A1 (\counter[0] ), .A2 (n_0_350), .B1 (n_0_440), .B2 (n_0_349));
AOI22_X1 i_0_516 (.ZN (n_0_324), .A1 (hfn_ipo_n79), .A2 (n_0_352), .B1 (hfn_ipo_n94), .B2 (n_0_351));
AOI22_X1 i_0_515 (.ZN (n_0_323), .A1 (hfn_ipo_n79), .A2 (n_0_348), .B1 (hfn_ipo_n94), .B2 (n_0_347));
AOI221_X1 i_0_514 (.ZN (n_0_322), .A (hfn_ipo_n65), .B1 (hfn_ipo_n71), .B2 (n_0_323)
    , .C1 (hfn_ipo_n69), .C2 (n_0_325));
AOI221_X1 i_0_513 (.ZN (n_0_321), .A (hfn_ipo_n67), .B1 (hfn_ipo_n71), .B2 (n_0_324)
    , .C1 (hfn_ipo_n69), .C2 (n_0_326));
NOR3_X1 i_0_512 (.ZN (n_0_320), .A1 (n_0_322), .A2 (n_0_321), .A3 (hfn_ipo_n75));
AOI221_X1 i_0_511 (.ZN (n_0_319), .A (hfn_ipo_n69), .B1 (hfn_ipo_n94), .B2 (n_0_355)
    , .C1 (hfn_ipo_n79), .C2 (n_0_356));
AOI221_X1 i_0_510 (.ZN (n_0_318), .A (hfn_ipo_n71), .B1 (\counter[0] ), .B2 (n_0_358)
    , .C1 (n_0_440), .C2 (n_0_357));
AOI221_X1 i_0_509 (.ZN (n_0_317), .A (hfn_ipo_n69), .B1 (hfn_ipo_n94), .B2 (n_0_359)
    , .C1 (hfn_ipo_n79), .C2 (n_0_360));
AOI221_X1 i_0_508 (.ZN (n_0_316), .A (hfn_ipo_n71), .B1 (\counter[0] ), .B2 (n_0_362)
    , .C1 (hfn_ipo_n94), .C2 (n_0_361));
OAI33_X1 i_0_507 (.ZN (n_0_315), .A1 (n_0_319), .A2 (n_0_318), .A3 (hfn_ipo_n65), .B1 (hfn_ipo_n67)
    , .B2 (n_0_316), .B3 (n_0_317));
NOR2_X1 i_0_506 (.ZN (n_0_314), .A1 (hfn_ipo_n77), .A2 (n_0_315));
AOI221_X1 i_0_505 (.ZN (n_0_313), .A (hfn_ipo_n71), .B1 (n_0_440), .B2 (n_0_345), .C1 (\counter[0] ), .C2 (n_0_346));
AOI221_X1 i_0_504 (.ZN (n_0_312), .A (hfn_ipo_n69), .B1 (hfn_ipo_n94), .B2 (n_0_343)
    , .C1 (hfn_ipo_n79), .C2 (n_0_344));
NOR3_X1 i_0_503 (.ZN (n_0_311), .A1 (hfn_ipo_n67), .A2 (n_0_312), .A3 (n_0_313));
AOI221_X1 i_0_502 (.ZN (n_0_310), .A (hfn_ipo_n69), .B1 (hfn_ipo_n94), .B2 (n_0_339)
    , .C1 (hfn_ipo_n79), .C2 (n_0_340));
AOI221_X1 i_0_501 (.ZN (n_0_309), .A (hfn_ipo_n71), .B1 (hfn_ipo_n94), .B2 (n_0_341)
    , .C1 (\counter[0] ), .C2 (n_0_342));
NOR3_X1 i_0_500 (.ZN (n_0_308), .A1 (hfn_ipo_n65), .A2 (n_0_309), .A3 (n_0_310));
NOR3_X1 i_0_499 (.ZN (n_0_307), .A1 (hfn_ipo_n77), .A2 (n_0_308), .A3 (n_0_311));
AOI22_X1 i_0_498 (.ZN (n_0_306), .A1 (\counter[0] ), .A2 (n_0_338), .B1 (n_0_440), .B2 (n_0_337));
OAI221_X1 i_0_497 (.ZN (n_0_305), .A (hfn_ipo_n71), .B1 (hfn_ipo_n94), .B2 (n_327)
    , .C1 (hfn_ipo_n79), .C2 (n_326));
AOI21_X1 i_0_496 (.ZN (n_0_304), .A (hfn_ipo_n67), .B1 (hfn_ipo_n69), .B2 (n_0_306));
AOI22_X1 i_0_495 (.ZN (n_0_303), .A1 (n_0_440), .A2 (n_0_333), .B1 (\counter[0] ), .B2 (n_0_334));
AOI22_X1 i_0_494 (.ZN (n_0_302), .A1 (hfn_ipo_n79), .A2 (n_0_332), .B1 (hfn_ipo_n94), .B2 (n_0_331));
AOI221_X1 i_0_493 (.ZN (n_0_301), .A (hfn_ipo_n65), .B1 (hfn_ipo_n71), .B2 (n_0_302)
    , .C1 (hfn_ipo_n69), .C2 (n_0_303));
AOI211_X1 i_0_492 (.ZN (n_0_300), .A (hfn_ipo_n75), .B (n_0_301), .C1 (n_0_305), .C2 (n_0_304));
OAI33_X1 i_0_491 (.ZN (n_0_299), .A1 (n_0_320), .A2 (n_0_314), .A3 (hfn_ipo_n83), .B1 (n_0_307)
    , .B2 (n_0_300), .B3 (hfn_ipo_n81));
INV_X1 i_0_490 (.ZN (n_0_298), .A (drc_ipo_n96));
AOI221_X1 i_0_489 (.ZN (n_0_297), .A (hfn_ipo_n76), .B1 (n_0_433), .B2 (n_0_369), .C1 (n_0_417), .C2 (hfn_ipo_n82));
OAI22_X1 i_0_488 (.ZN (n_0_296), .A1 (n_0_409), .A2 (hfn_ipo_n83), .B1 (n_0_425), .B2 (hfn_ipo_n82));
AOI21_X1 i_0_487 (.ZN (n_0_295), .A (n_0_297), .B1 (hfn_ipo_n76), .B2 (n_0_296));
OAI22_X1 i_0_486 (.ZN (n_0_294), .A1 (n_0_405), .A2 (hfn_ipo_n83), .B1 (n_0_421), .B2 (hfn_ipo_n82));
AOI221_X1 i_0_485 (.ZN (n_0_293), .A (hfn_ipo_n76), .B1 (n_0_413), .B2 (hfn_ipo_n82)
    , .C1 (n_0_429), .C2 (n_0_369));
AOI21_X1 i_0_484 (.ZN (n_0_292), .A (n_0_293), .B1 (hfn_ipo_n76), .B2 (n_0_294));
AOI221_X1 i_0_483 (.ZN (n_0_291), .A (hfn_ipo_n70), .B1 (hfn_ipo_n66), .B2 (n_0_292)
    , .C1 (hfn_ipo_n68), .C2 (n_0_295));
AOI221_X1 i_0_482 (.ZN (n_0_290), .A (hfn_ipo_n76), .B1 (n_0_431), .B2 (n_0_369), .C1 (n_0_415), .C2 (hfn_ipo_n82));
OAI22_X1 i_0_481 (.ZN (n_0_289), .A1 (n_0_407), .A2 (n_0_369), .B1 (n_0_423), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_480 (.ZN (n_0_288), .A1 (n_0_403), .A2 (n_0_369), .B1 (n_0_419), .B2 (hfn_ipo_n82));
AOI221_X1 i_0_479 (.ZN (n_0_287), .A (hfn_ipo_n76), .B1 (n_0_411), .B2 (hfn_ipo_n82)
    , .C1 (n_0_427), .C2 (n_0_369));
AOI21_X1 i_0_478 (.ZN (n_0_286), .A (n_0_287), .B1 (hfn_ipo_n76), .B2 (n_0_288));
AOI211_X1 i_0_477 (.ZN (n_0_285), .A (n_0_290), .B (hfn_ipo_n66), .C1 (hfn_ipo_n76), .C2 (n_0_289));
AOI21_X1 i_0_476 (.ZN (n_0_284), .A (n_0_285), .B1 (hfn_ipo_n66), .B2 (n_0_286));
OAI22_X1 i_0_475 (.ZN (n_0_283), .A1 (n_0_408), .A2 (n_0_369), .B1 (n_0_424), .B2 (hfn_ipo_n82));
AOI221_X1 i_0_474 (.ZN (n_0_282), .A (hfn_ipo_n76), .B1 (n_0_416), .B2 (hfn_ipo_n82)
    , .C1 (n_0_432), .C2 (n_0_369));
AOI211_X1 i_0_473 (.ZN (n_0_281), .A (hfn_ipo_n66), .B (n_0_282), .C1 (hfn_ipo_n76), .C2 (n_0_283));
OAI22_X1 i_0_472 (.ZN (n_0_280), .A1 (n_0_404), .A2 (n_0_369), .B1 (n_0_420), .B2 (hfn_ipo_n82));
AOI221_X1 i_0_471 (.ZN (n_0_279), .A (hfn_ipo_n76), .B1 (n_0_412), .B2 (hfn_ipo_n82)
    , .C1 (n_0_428), .C2 (n_0_369));
AOI21_X1 i_0_470 (.ZN (n_0_278), .A (n_0_279), .B1 (hfn_ipo_n76), .B2 (n_0_280));
AOI221_X1 i_0_469 (.ZN (n_0_277), .A (hfn_ipo_n75), .B1 (n_0_414), .B2 (hfn_ipo_n82)
    , .C1 (n_0_430), .C2 (n_0_369));
OAI22_X1 i_0_468 (.ZN (n_0_276), .A1 (n_0_406), .A2 (hfn_ipo_n83), .B1 (n_0_422), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_467 (.ZN (n_0_275), .A1 (n_0_402), .A2 (hfn_ipo_n83), .B1 (n_0_418), .B2 (hfn_ipo_n81));
AOI221_X1 i_0_466 (.ZN (n_0_274), .A (hfn_ipo_n76), .B1 (n_0_410), .B2 (hfn_ipo_n82)
    , .C1 (n_0_426), .C2 (n_0_369));
AOI21_X1 i_0_465 (.ZN (n_0_273), .A (n_0_274), .B1 (hfn_ipo_n76), .B2 (n_0_275));
AOI211_X1 i_0_464 (.ZN (n_0_272), .A (n_0_277), .B (hfn_ipo_n66), .C1 (hfn_ipo_n75), .C2 (n_0_276));
AOI21_X1 i_0_463 (.ZN (n_0_271), .A (n_0_272), .B1 (hfn_ipo_n66), .B2 (n_0_273));
AOI211_X1 i_0_462 (.ZN (n_0_270), .A (n_0_281), .B (hfn_ipo_n70), .C1 (hfn_ipo_n66), .C2 (n_0_278));
AOI21_X1 i_0_461 (.ZN (n_0_269), .A (n_0_270), .B1 (hfn_ipo_n70), .B2 (n_0_271));
AOI211_X1 i_0_460 (.ZN (n_0_268), .A (n_0_291), .B (hfn_ipo_n80), .C1 (hfn_ipo_n70), .C2 (n_0_284));
AOI211_X1 i_0_459 (.ZN (n_321), .A (n_0_268), .B (drc_ipo_n96), .C1 (hfn_ipo_n80), .C2 (n_0_269));
OAI22_X1 i_0_458 (.ZN (n_0_267), .A1 (n_0_401), .A2 (n_0_369), .B1 (n_0_417), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_457 (.ZN (n_0_266), .A1 (hfn_ipo_n76), .A2 (n_0_267), .B1 (hfn_ipo_n78), .B2 (n_0_296));
OAI22_X1 i_0_456 (.ZN (n_0_265), .A1 (hfn_ipo_n66), .A2 (n_0_292), .B1 (hfn_ipo_n68), .B2 (n_0_266));
AOI22_X1 i_0_455 (.ZN (n_0_264), .A1 (hfn_ipo_n72), .A2 (n_0_284), .B1 (hfn_ipo_n70), .B2 (n_0_265));
AOI221_X1 i_0_454 (.ZN (n_320), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_264)
    , .C1 (hfn_ipo_n95), .C2 (n_0_269));
OAI22_X1 i_0_453 (.ZN (n_0_263), .A1 (n_0_416), .A2 (hfn_ipo_n82), .B1 (n_0_400), .B2 (n_0_369));
AOI22_X1 i_0_452 (.ZN (n_0_262), .A1 (hfn_ipo_n76), .A2 (n_0_263), .B1 (hfn_ipo_n78), .B2 (n_0_283));
OAI22_X1 i_0_451 (.ZN (n_0_261), .A1 (hfn_ipo_n66), .A2 (n_0_278), .B1 (hfn_ipo_n68), .B2 (n_0_262));
AOI22_X1 i_0_450 (.ZN (n_0_260), .A1 (hfn_ipo_n72), .A2 (n_0_271), .B1 (hfn_ipo_n70), .B2 (n_0_261));
AOI221_X1 i_0_449 (.ZN (n_319), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_264)
    , .C1 (hfn_ipo_n80), .C2 (n_0_260));
OAI22_X1 i_0_448 (.ZN (n_0_259), .A1 (n_0_415), .A2 (hfn_ipo_n82), .B1 (n_0_399), .B2 (n_0_369));
AOI22_X1 i_0_447 (.ZN (n_0_258), .A1 (hfn_ipo_n76), .A2 (n_0_259), .B1 (hfn_ipo_n78), .B2 (n_0_289));
OAI22_X1 i_0_446 (.ZN (n_0_257), .A1 (hfn_ipo_n66), .A2 (n_0_286), .B1 (hfn_ipo_n68), .B2 (n_0_258));
AOI22_X1 i_0_445 (.ZN (n_0_256), .A1 (hfn_ipo_n72), .A2 (n_0_265), .B1 (hfn_ipo_n70), .B2 (n_0_257));
AOI221_X1 i_0_444 (.ZN (n_318), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_260)
    , .C1 (hfn_ipo_n80), .C2 (n_0_256));
OAI22_X1 i_0_443 (.ZN (n_0_255), .A1 (n_0_414), .A2 (hfn_ipo_n82), .B1 (n_0_398), .B2 (n_0_369));
AOI22_X1 i_0_442 (.ZN (n_0_254), .A1 (hfn_ipo_n76), .A2 (n_0_255), .B1 (hfn_ipo_n78), .B2 (n_0_276));
OAI22_X1 i_0_441 (.ZN (n_0_253), .A1 (hfn_ipo_n66), .A2 (n_0_273), .B1 (hfn_ipo_n68), .B2 (n_0_254));
AOI22_X1 i_0_440 (.ZN (n_0_252), .A1 (hfn_ipo_n70), .A2 (n_0_253), .B1 (hfn_ipo_n72), .B2 (n_0_261));
AOI221_X1 i_0_439 (.ZN (n_317), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_256)
    , .C1 (hfn_ipo_n80), .C2 (n_0_252));
OAI22_X1 i_0_438 (.ZN (n_0_251), .A1 (n_0_413), .A2 (hfn_ipo_n82), .B1 (n_0_397), .B2 (n_0_369));
AOI22_X1 i_0_437 (.ZN (n_0_250), .A1 (hfn_ipo_n76), .A2 (n_0_251), .B1 (hfn_ipo_n78), .B2 (n_0_294));
OAI22_X1 i_0_436 (.ZN (n_0_249), .A1 (hfn_ipo_n66), .A2 (n_0_266), .B1 (hfn_ipo_n68), .B2 (n_0_250));
AOI22_X1 i_0_435 (.ZN (n_0_248), .A1 (hfn_ipo_n72), .A2 (n_0_257), .B1 (hfn_ipo_n70), .B2 (n_0_249));
AOI221_X1 i_0_434 (.ZN (n_316), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_252)
    , .C1 (hfn_ipo_n80), .C2 (n_0_248));
OAI22_X1 i_0_433 (.ZN (n_0_247), .A1 (n_0_412), .A2 (hfn_ipo_n82), .B1 (n_0_396), .B2 (n_0_369));
AOI22_X1 i_0_432 (.ZN (n_0_246), .A1 (hfn_ipo_n76), .A2 (n_0_247), .B1 (hfn_ipo_n78), .B2 (n_0_280));
OAI22_X1 i_0_431 (.ZN (n_0_245), .A1 (hfn_ipo_n68), .A2 (n_0_246), .B1 (hfn_ipo_n66), .B2 (n_0_262));
AOI22_X1 i_0_430 (.ZN (n_0_244), .A1 (hfn_ipo_n72), .A2 (n_0_253), .B1 (hfn_ipo_n70), .B2 (n_0_245));
AOI221_X1 i_0_429 (.ZN (n_315), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_244)
    , .C1 (hfn_ipo_n95), .C2 (n_0_248));
OAI22_X1 i_0_428 (.ZN (n_0_243), .A1 (n_0_411), .A2 (hfn_ipo_n82), .B1 (n_0_395), .B2 (n_0_369));
AOI22_X1 i_0_427 (.ZN (n_0_242), .A1 (hfn_ipo_n76), .A2 (n_0_243), .B1 (hfn_ipo_n78), .B2 (n_0_288));
OAI22_X1 i_0_426 (.ZN (n_0_241), .A1 (hfn_ipo_n68), .A2 (n_0_242), .B1 (hfn_ipo_n66), .B2 (n_0_258));
AOI22_X1 i_0_425 (.ZN (n_0_240), .A1 (hfn_ipo_n72), .A2 (n_0_249), .B1 (hfn_ipo_n70), .B2 (n_0_241));
AOI221_X1 i_0_424 (.ZN (n_314), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_240)
    , .C1 (hfn_ipo_n95), .C2 (n_0_244));
OAI22_X1 i_0_423 (.ZN (n_0_239), .A1 (n_0_410), .A2 (hfn_ipo_n82), .B1 (n_0_394), .B2 (n_0_369));
AOI22_X1 i_0_422 (.ZN (n_0_238), .A1 (hfn_ipo_n75), .A2 (n_0_239), .B1 (hfn_ipo_n78), .B2 (n_0_275));
OAI22_X1 i_0_421 (.ZN (n_0_237), .A1 (hfn_ipo_n68), .A2 (n_0_238), .B1 (hfn_ipo_n66), .B2 (n_0_254));
AOI22_X1 i_0_420 (.ZN (n_0_236), .A1 (hfn_ipo_n70), .A2 (n_0_237), .B1 (hfn_ipo_n72), .B2 (n_0_245));
AOI221_X1 i_0_419 (.ZN (n_313), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_236)
    , .C1 (hfn_ipo_n95), .C2 (n_0_240));
OAI22_X1 i_0_418 (.ZN (n_0_235), .A1 (n_0_409), .A2 (hfn_ipo_n81), .B1 (n_0_393), .B2 (hfn_ipo_n83));
AOI22_X1 i_0_417 (.ZN (n_0_234), .A1 (hfn_ipo_n78), .A2 (n_0_267), .B1 (hfn_ipo_n76), .B2 (n_0_235));
OAI22_X1 i_0_416 (.ZN (n_0_233), .A1 (hfn_ipo_n66), .A2 (n_0_250), .B1 (hfn_ipo_n68), .B2 (n_0_234));
AOI22_X1 i_0_415 (.ZN (n_0_232), .A1 (hfn_ipo_n70), .A2 (n_0_233), .B1 (hfn_ipo_n72), .B2 (n_0_241));
AOI221_X1 i_0_414 (.ZN (n_312), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_236)
    , .C1 (hfn_ipo_n80), .C2 (n_0_232));
OAI22_X1 i_0_413 (.ZN (n_0_231), .A1 (n_0_408), .A2 (hfn_ipo_n82), .B1 (n_0_392), .B2 (n_0_369));
AOI22_X1 i_0_412 (.ZN (n_0_230), .A1 (hfn_ipo_n76), .A2 (n_0_231), .B1 (hfn_ipo_n78), .B2 (n_0_263));
OAI22_X1 i_0_411 (.ZN (n_0_229), .A1 (hfn_ipo_n66), .A2 (n_0_246), .B1 (hfn_ipo_n68), .B2 (n_0_230));
AOI22_X1 i_0_410 (.ZN (n_0_228), .A1 (hfn_ipo_n70), .A2 (n_0_229), .B1 (hfn_ipo_n72), .B2 (n_0_237));
AOI221_X1 i_0_409 (.ZN (n_311), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_232)
    , .C1 (hfn_ipo_n80), .C2 (n_0_228));
OAI22_X1 i_0_408 (.ZN (n_0_227), .A1 (n_0_407), .A2 (hfn_ipo_n82), .B1 (n_0_391), .B2 (n_0_369));
AOI22_X1 i_0_407 (.ZN (n_0_226), .A1 (hfn_ipo_n76), .A2 (n_0_227), .B1 (hfn_ipo_n78), .B2 (n_0_259));
OAI22_X1 i_0_406 (.ZN (n_0_225), .A1 (hfn_ipo_n66), .A2 (n_0_242), .B1 (hfn_ipo_n68), .B2 (n_0_226));
AOI22_X1 i_0_405 (.ZN (n_0_224), .A1 (hfn_ipo_n72), .A2 (n_0_233), .B1 (hfn_ipo_n70), .B2 (n_0_225));
AOI221_X1 i_0_404 (.ZN (n_310), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_228)
    , .C1 (hfn_ipo_n80), .C2 (n_0_224));
OAI22_X1 i_0_403 (.ZN (n_0_223), .A1 (n_0_406), .A2 (hfn_ipo_n81), .B1 (n_0_390), .B2 (hfn_ipo_n83));
AOI22_X1 i_0_402 (.ZN (n_0_222), .A1 (hfn_ipo_n76), .A2 (n_0_223), .B1 (hfn_ipo_n78), .B2 (n_0_255));
OAI22_X1 i_0_401 (.ZN (n_0_221), .A1 (hfn_ipo_n66), .A2 (n_0_238), .B1 (hfn_ipo_n68), .B2 (n_0_222));
AOI22_X1 i_0_400 (.ZN (n_0_220), .A1 (hfn_ipo_n70), .A2 (n_0_221), .B1 (hfn_ipo_n72), .B2 (n_0_229));
AOI221_X1 i_0_399 (.ZN (n_309), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_224)
    , .C1 (hfn_ipo_n80), .C2 (n_0_220));
OAI22_X1 i_0_398 (.ZN (n_0_219), .A1 (n_0_405), .A2 (hfn_ipo_n82), .B1 (n_0_389), .B2 (hfn_ipo_n83));
AOI22_X1 i_0_397 (.ZN (n_0_218), .A1 (hfn_ipo_n76), .A2 (n_0_219), .B1 (hfn_ipo_n78), .B2 (n_0_251));
OAI22_X1 i_0_396 (.ZN (n_0_217), .A1 (hfn_ipo_n66), .A2 (n_0_234), .B1 (hfn_ipo_n68), .B2 (n_0_218));
AOI22_X1 i_0_395 (.ZN (n_0_216), .A1 (hfn_ipo_n70), .A2 (n_0_217), .B1 (hfn_ipo_n72), .B2 (n_0_225));
AOI221_X1 i_0_394 (.ZN (n_308), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_220)
    , .C1 (hfn_ipo_n80), .C2 (n_0_216));
OAI22_X1 i_0_393 (.ZN (n_0_215), .A1 (n_0_404), .A2 (hfn_ipo_n82), .B1 (n_0_388), .B2 (n_0_369));
AOI22_X1 i_0_392 (.ZN (n_0_214), .A1 (hfn_ipo_n76), .A2 (n_0_215), .B1 (hfn_ipo_n78), .B2 (n_0_247));
OAI22_X1 i_0_391 (.ZN (n_0_213), .A1 (hfn_ipo_n68), .A2 (n_0_214), .B1 (hfn_ipo_n66), .B2 (n_0_230));
AOI22_X1 i_0_390 (.ZN (n_0_212), .A1 (hfn_ipo_n72), .A2 (n_0_221), .B1 (hfn_ipo_n70), .B2 (n_0_213));
AOI221_X1 i_0_389 (.ZN (n_307), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_212)
    , .C1 (hfn_ipo_n95), .C2 (n_0_216));
OAI22_X1 i_0_388 (.ZN (n_0_211), .A1 (n_0_403), .A2 (hfn_ipo_n82), .B1 (n_0_387), .B2 (n_0_369));
AOI22_X1 i_0_387 (.ZN (n_0_210), .A1 (hfn_ipo_n76), .A2 (n_0_211), .B1 (hfn_ipo_n78), .B2 (n_0_243));
OAI22_X1 i_0_386 (.ZN (n_0_209), .A1 (hfn_ipo_n68), .A2 (n_0_210), .B1 (hfn_ipo_n66), .B2 (n_0_226));
AOI22_X1 i_0_385 (.ZN (n_0_208), .A1 (hfn_ipo_n72), .A2 (n_0_217), .B1 (hfn_ipo_n70), .B2 (n_0_209));
AOI221_X1 i_0_384 (.ZN (n_306), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_212)
    , .C1 (hfn_ipo_n80), .C2 (n_0_208));
OAI22_X1 i_0_383 (.ZN (n_0_207), .A1 (n_0_402), .A2 (hfn_ipo_n81), .B1 (n_0_386), .B2 (hfn_ipo_n83));
AOI22_X1 i_0_382 (.ZN (n_0_206), .A1 (hfn_ipo_n75), .A2 (n_0_207), .B1 (hfn_ipo_n78), .B2 (n_0_239));
OAI22_X1 i_0_381 (.ZN (n_0_205), .A1 (hfn_ipo_n68), .A2 (n_0_206), .B1 (hfn_ipo_n66), .B2 (n_0_222));
AOI22_X1 i_0_380 (.ZN (n_0_204), .A1 (hfn_ipo_n70), .A2 (n_0_205), .B1 (hfn_ipo_n72), .B2 (n_0_213));
AOI221_X1 i_0_379 (.ZN (n_305), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_204)
    , .C1 (hfn_ipo_n95), .C2 (n_0_208));
OAI22_X1 i_0_378 (.ZN (n_0_203), .A1 (n_0_401), .A2 (hfn_ipo_n82), .B1 (n_0_385), .B2 (hfn_ipo_n83));
AOI22_X1 i_0_377 (.ZN (n_0_202), .A1 (hfn_ipo_n76), .A2 (n_0_203), .B1 (hfn_ipo_n78), .B2 (n_0_235));
OAI22_X1 i_0_376 (.ZN (n_0_201), .A1 (hfn_ipo_n68), .A2 (n_0_202), .B1 (hfn_ipo_n66), .B2 (n_0_218));
AOI22_X1 i_0_375 (.ZN (n_0_200), .A1 (hfn_ipo_n70), .A2 (n_0_201), .B1 (hfn_ipo_n72), .B2 (n_0_209));
AOI221_X1 i_0_374 (.ZN (n_304), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_204)
    , .C1 (hfn_ipo_n80), .C2 (n_0_200));
OAI22_X1 i_0_373 (.ZN (n_0_199), .A1 (n_0_384), .A2 (n_0_369), .B1 (n_0_400), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_372 (.ZN (n_0_198), .A1 (hfn_ipo_n78), .A2 (n_0_231), .B1 (hfn_ipo_n76), .B2 (n_0_199));
OAI22_X1 i_0_371 (.ZN (n_0_197), .A1 (hfn_ipo_n66), .A2 (n_0_214), .B1 (hfn_ipo_n68), .B2 (n_0_198));
AOI22_X1 i_0_370 (.ZN (n_0_196), .A1 (hfn_ipo_n72), .A2 (n_0_205), .B1 (hfn_ipo_n70), .B2 (n_0_197));
AOI221_X1 i_0_369 (.ZN (n_303), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_200)
    , .C1 (hfn_ipo_n80), .C2 (n_0_196));
OAI22_X1 i_0_368 (.ZN (n_0_195), .A1 (n_0_383), .A2 (n_0_369), .B1 (n_0_399), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_367 (.ZN (n_0_194), .A1 (hfn_ipo_n78), .A2 (n_0_227), .B1 (hfn_ipo_n76), .B2 (n_0_195));
OAI22_X1 i_0_366 (.ZN (n_0_193), .A1 (hfn_ipo_n66), .A2 (n_0_210), .B1 (hfn_ipo_n68), .B2 (n_0_194));
AOI22_X1 i_0_365 (.ZN (n_0_192), .A1 (hfn_ipo_n72), .A2 (n_0_201), .B1 (hfn_ipo_n70), .B2 (n_0_193));
AOI221_X1 i_0_364 (.ZN (n_302), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_196)
    , .C1 (hfn_ipo_n80), .C2 (n_0_192));
OAI22_X1 i_0_363 (.ZN (n_0_191), .A1 (n_0_382), .A2 (hfn_ipo_n83), .B1 (n_0_398), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_362 (.ZN (n_0_190), .A1 (hfn_ipo_n78), .A2 (n_0_223), .B1 (hfn_ipo_n75), .B2 (n_0_191));
OAI22_X1 i_0_361 (.ZN (n_0_189), .A1 (hfn_ipo_n66), .A2 (n_0_206), .B1 (hfn_ipo_n68), .B2 (n_0_190));
AOI22_X1 i_0_360 (.ZN (n_0_188), .A1 (hfn_ipo_n70), .A2 (n_0_189), .B1 (hfn_ipo_n72), .B2 (n_0_197));
AOI221_X1 i_0_359 (.ZN (n_301), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_192)
    , .C1 (hfn_ipo_n80), .C2 (n_0_188));
OAI22_X1 i_0_358 (.ZN (n_0_187), .A1 (n_0_381), .A2 (hfn_ipo_n83), .B1 (n_0_397), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_357 (.ZN (n_0_186), .A1 (hfn_ipo_n78), .A2 (n_0_219), .B1 (hfn_ipo_n75), .B2 (n_0_187));
OAI22_X1 i_0_356 (.ZN (n_0_185), .A1 (hfn_ipo_n66), .A2 (n_0_202), .B1 (hfn_ipo_n68), .B2 (n_0_186));
AOI22_X1 i_0_355 (.ZN (n_0_184), .A1 (hfn_ipo_n70), .A2 (n_0_185), .B1 (hfn_ipo_n72), .B2 (n_0_193));
AOI221_X1 i_0_354 (.ZN (n_300), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_188)
    , .C1 (hfn_ipo_n80), .C2 (n_0_184));
OAI22_X1 i_0_353 (.ZN (n_0_183), .A1 (n_0_380), .A2 (hfn_ipo_n83), .B1 (n_0_396), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_352 (.ZN (n_0_182), .A1 (hfn_ipo_n78), .A2 (n_0_215), .B1 (hfn_ipo_n76), .B2 (n_0_183));
OAI22_X1 i_0_351 (.ZN (n_0_181), .A1 (hfn_ipo_n68), .A2 (n_0_182), .B1 (hfn_ipo_n66), .B2 (n_0_198));
AOI22_X1 i_0_350 (.ZN (n_0_180), .A1 (hfn_ipo_n70), .A2 (n_0_181), .B1 (hfn_ipo_n72), .B2 (n_0_189));
AOI221_X1 i_0_349 (.ZN (n_299), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_180)
    , .C1 (hfn_ipo_n95), .C2 (n_0_184));
OAI22_X1 i_0_348 (.ZN (n_0_179), .A1 (n_0_379), .A2 (hfn_ipo_n83), .B1 (n_0_395), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_347 (.ZN (n_0_178), .A1 (hfn_ipo_n78), .A2 (n_0_211), .B1 (hfn_ipo_n76), .B2 (n_0_179));
OAI22_X1 i_0_346 (.ZN (n_0_177), .A1 (hfn_ipo_n68), .A2 (n_0_178), .B1 (hfn_ipo_n66), .B2 (n_0_194));
AOI22_X1 i_0_345 (.ZN (n_0_176), .A1 (hfn_ipo_n72), .A2 (n_0_185), .B1 (hfn_ipo_n70), .B2 (n_0_177));
AOI221_X1 i_0_344 (.ZN (n_298), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_176)
    , .C1 (hfn_ipo_n95), .C2 (n_0_180));
OAI22_X1 i_0_343 (.ZN (n_0_175), .A1 (n_0_378), .A2 (hfn_ipo_n83), .B1 (n_0_394), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_342 (.ZN (n_0_174), .A1 (hfn_ipo_n78), .A2 (n_0_207), .B1 (hfn_ipo_n75), .B2 (n_0_175));
OAI22_X1 i_0_341 (.ZN (n_0_173), .A1 (hfn_ipo_n68), .A2 (n_0_174), .B1 (hfn_ipo_n66), .B2 (n_0_190));
AOI22_X1 i_0_340 (.ZN (n_0_172), .A1 (hfn_ipo_n70), .A2 (n_0_173), .B1 (hfn_ipo_n72), .B2 (n_0_181));
AOI221_X1 i_0_339 (.ZN (n_297), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_172)
    , .C1 (hfn_ipo_n95), .C2 (n_0_176));
OAI22_X1 i_0_338 (.ZN (n_0_171), .A1 (n_0_377), .A2 (hfn_ipo_n83), .B1 (n_0_393), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_337 (.ZN (n_0_170), .A1 (hfn_ipo_n78), .A2 (n_0_203), .B1 (hfn_ipo_n75), .B2 (n_0_171));
OAI22_X1 i_0_336 (.ZN (n_0_169), .A1 (hfn_ipo_n68), .A2 (n_0_170), .B1 (hfn_ipo_n66), .B2 (n_0_186));
AOI22_X1 i_0_335 (.ZN (n_0_168), .A1 (hfn_ipo_n70), .A2 (n_0_169), .B1 (hfn_ipo_n72), .B2 (n_0_177));
AOI221_X1 i_0_334 (.ZN (n_296), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_168)
    , .C1 (hfn_ipo_n95), .C2 (n_0_172));
OAI22_X1 i_0_333 (.ZN (n_0_167), .A1 (n_0_376), .A2 (hfn_ipo_n83), .B1 (n_0_392), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_332 (.ZN (n_0_166), .A1 (hfn_ipo_n75), .A2 (n_0_167), .B1 (hfn_ipo_n78), .B2 (n_0_199));
OAI22_X1 i_0_331 (.ZN (n_0_165), .A1 (hfn_ipo_n68), .A2 (n_0_166), .B1 (hfn_ipo_n66), .B2 (n_0_182));
AOI22_X1 i_0_330 (.ZN (n_0_164), .A1 (hfn_ipo_n70), .A2 (n_0_165), .B1 (hfn_ipo_n72), .B2 (n_0_173));
AOI221_X1 i_0_329 (.ZN (n_295), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_168)
    , .C1 (hfn_ipo_n80), .C2 (n_0_164));
OAI22_X1 i_0_328 (.ZN (n_0_163), .A1 (n_0_375), .A2 (hfn_ipo_n83), .B1 (n_0_391), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_327 (.ZN (n_0_162), .A1 (hfn_ipo_n75), .A2 (n_0_163), .B1 (hfn_ipo_n78), .B2 (n_0_195));
OAI22_X1 i_0_326 (.ZN (n_0_161), .A1 (hfn_ipo_n68), .A2 (n_0_162), .B1 (hfn_ipo_n66), .B2 (n_0_178));
AOI22_X1 i_0_325 (.ZN (n_0_160), .A1 (hfn_ipo_n72), .A2 (n_0_169), .B1 (hfn_ipo_n70), .B2 (n_0_161));
AOI221_X1 i_0_324 (.ZN (n_294), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_160)
    , .C1 (hfn_ipo_n95), .C2 (n_0_164));
OAI22_X1 i_0_323 (.ZN (n_0_159), .A1 (n_0_374), .A2 (hfn_ipo_n83), .B1 (n_0_390), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_322 (.ZN (n_0_158), .A1 (hfn_ipo_n75), .A2 (n_0_159), .B1 (hfn_ipo_n78), .B2 (n_0_191));
OAI22_X1 i_0_321 (.ZN (n_0_157), .A1 (hfn_ipo_n68), .A2 (n_0_158), .B1 (hfn_ipo_n66), .B2 (n_0_174));
AOI22_X1 i_0_320 (.ZN (n_0_156), .A1 (hfn_ipo_n70), .A2 (n_0_157), .B1 (hfn_ipo_n72), .B2 (n_0_165));
AOI221_X1 i_0_319 (.ZN (n_293), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_160)
    , .C1 (hfn_ipo_n80), .C2 (n_0_156));
OAI22_X1 i_0_318 (.ZN (n_0_155), .A1 (n_0_373), .A2 (hfn_ipo_n83), .B1 (n_0_389), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_317 (.ZN (n_0_154), .A1 (hfn_ipo_n75), .A2 (n_0_155), .B1 (hfn_ipo_n78), .B2 (n_0_187));
OAI22_X1 i_0_316 (.ZN (n_0_153), .A1 (hfn_ipo_n65), .A2 (n_0_170), .B1 (hfn_ipo_n67), .B2 (n_0_154));
AOI22_X1 i_0_315 (.ZN (n_0_152), .A1 (hfn_ipo_n70), .A2 (n_0_153), .B1 (hfn_ipo_n72), .B2 (n_0_161));
AOI221_X1 i_0_314 (.ZN (n_292), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_156)
    , .C1 (hfn_ipo_n80), .C2 (n_0_152));
OAI22_X1 i_0_313 (.ZN (n_0_151), .A1 (n_0_372), .A2 (hfn_ipo_n83), .B1 (n_0_388), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_312 (.ZN (n_0_150), .A1 (hfn_ipo_n75), .A2 (n_0_151), .B1 (hfn_ipo_n78), .B2 (n_0_183));
OAI22_X1 i_0_311 (.ZN (n_0_149), .A1 (hfn_ipo_n68), .A2 (n_0_150), .B1 (hfn_ipo_n66), .B2 (n_0_166));
AOI22_X1 i_0_310 (.ZN (n_0_148), .A1 (hfn_ipo_n70), .A2 (n_0_149), .B1 (hfn_ipo_n72), .B2 (n_0_157));
AOI221_X1 i_0_309 (.ZN (n_291), .A (drc_ipo_n96), .B1 (hfn_ipo_n95), .B2 (n_0_152)
    , .C1 (hfn_ipo_n80), .C2 (n_0_148));
OAI22_X1 i_0_308 (.ZN (n_0_147), .A1 (n_0_371), .A2 (hfn_ipo_n83), .B1 (n_0_387), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_307 (.ZN (n_0_146), .A1 (hfn_ipo_n75), .A2 (n_0_147), .B1 (hfn_ipo_n77), .B2 (n_0_179));
OAI22_X1 i_0_306 (.ZN (n_0_145), .A1 (hfn_ipo_n68), .A2 (n_0_146), .B1 (hfn_ipo_n65), .B2 (n_0_162));
AOI22_X1 i_0_305 (.ZN (n_0_144), .A1 (hfn_ipo_n72), .A2 (n_0_153), .B1 (hfn_ipo_n70), .B2 (n_0_145));
AOI221_X1 i_0_304 (.ZN (n_290), .A (drc_ipo_n96), .B1 (hfn_ipo_n80), .B2 (n_0_144)
    , .C1 (hfn_ipo_n95), .C2 (n_0_148));
AOI22_X1 i_0_303 (.ZN (n_0_143), .A1 (n_0_386), .A2 (hfn_ipo_n83), .B1 (n_0_439), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_302 (.ZN (n_0_142), .A1 (hfn_ipo_n77), .A2 (n_0_175), .B1 (hfn_ipo_n75), .B2 (n_0_143));
OAI22_X1 i_0_301 (.ZN (n_0_141), .A1 (hfn_ipo_n65), .A2 (n_0_158), .B1 (hfn_ipo_n67), .B2 (n_0_142));
AOI22_X1 i_0_300 (.ZN (n_0_140), .A1 (hfn_ipo_n72), .A2 (n_0_149), .B1 (hfn_ipo_n70), .B2 (n_0_141));
OAI22_X1 i_0_299 (.ZN (n_0_139), .A1 (hfn_ipo_n95), .A2 (n_0_140), .B1 (hfn_ipo_n80), .B2 (n_0_144));
AND2_X1 i_0_298 (.ZN (n_289), .A1 (n_0_298), .A2 (n_0_139));
NOR2_X1 i_0_297 (.ZN (n_0_138), .A1 (n_0_385), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_296 (.ZN (n_0_137), .A1 (hfn_ipo_n77), .A2 (n_0_171), .B1 (hfn_ipo_n75), .B2 (n_0_138));
OAI22_X1 i_0_295 (.ZN (n_0_136), .A1 (hfn_ipo_n65), .A2 (n_0_154), .B1 (hfn_ipo_n67), .B2 (n_0_137));
AOI22_X1 i_0_294 (.ZN (n_0_135), .A1 (hfn_ipo_n72), .A2 (n_0_145), .B1 (hfn_ipo_n69), .B2 (n_0_136));
OAI22_X1 i_0_293 (.ZN (n_0_134), .A1 (hfn_ipo_n95), .A2 (n_0_135), .B1 (hfn_ipo_n80), .B2 (n_0_140));
AND2_X1 i_0_292 (.ZN (n_288), .A1 (n_0_298), .A2 (n_0_134));
NOR2_X1 i_0_291 (.ZN (n_0_133), .A1 (n_0_384), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_290 (.ZN (n_0_132), .A1 (hfn_ipo_n77), .A2 (n_0_167), .B1 (hfn_ipo_n75), .B2 (n_0_133));
OAI22_X1 i_0_289 (.ZN (n_0_131), .A1 (hfn_ipo_n65), .A2 (n_0_150), .B1 (hfn_ipo_n67), .B2 (n_0_132));
AOI22_X1 i_0_288 (.ZN (n_0_130), .A1 (hfn_ipo_n72), .A2 (n_0_141), .B1 (hfn_ipo_n69), .B2 (n_0_131));
OAI22_X1 i_0_287 (.ZN (n_0_129), .A1 (hfn_ipo_n95), .A2 (n_0_130), .B1 (hfn_ipo_n80), .B2 (n_0_135));
AND2_X1 i_0_286 (.ZN (n_287), .A1 (n_0_298), .A2 (n_0_129));
NOR2_X1 i_0_285 (.ZN (n_0_128), .A1 (n_0_383), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_284 (.ZN (n_0_127), .A1 (hfn_ipo_n77), .A2 (n_0_163), .B1 (hfn_ipo_n75), .B2 (n_0_128));
OAI22_X1 i_0_283 (.ZN (n_0_126), .A1 (hfn_ipo_n65), .A2 (n_0_146), .B1 (hfn_ipo_n67), .B2 (n_0_127));
AOI22_X1 i_0_282 (.ZN (n_0_125), .A1 (hfn_ipo_n69), .A2 (n_0_126), .B1 (hfn_ipo_n71), .B2 (n_0_136));
OAI22_X1 i_0_281 (.ZN (n_0_124), .A1 (hfn_ipo_n95), .A2 (n_0_125), .B1 (hfn_ipo_n80), .B2 (n_0_130));
AND2_X1 i_0_280 (.ZN (n_286), .A1 (n_0_298), .A2 (n_0_124));
NOR2_X1 i_0_279 (.ZN (n_0_123), .A1 (n_0_382), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_278 (.ZN (n_0_122), .A1 (hfn_ipo_n77), .A2 (n_0_159), .B1 (hfn_ipo_n75), .B2 (n_0_123));
OAI22_X1 i_0_277 (.ZN (n_0_121), .A1 (hfn_ipo_n65), .A2 (n_0_142), .B1 (hfn_ipo_n67), .B2 (n_0_122));
AOI22_X1 i_0_276 (.ZN (n_0_120), .A1 (hfn_ipo_n71), .A2 (n_0_131), .B1 (hfn_ipo_n69), .B2 (n_0_121));
OAI22_X1 i_0_275 (.ZN (n_0_119), .A1 (hfn_ipo_n95), .A2 (n_0_120), .B1 (hfn_ipo_n79), .B2 (n_0_125));
AND2_X1 i_0_274 (.ZN (n_285), .A1 (n_0_298), .A2 (n_0_119));
NOR2_X1 i_0_273 (.ZN (n_0_118), .A1 (n_0_381), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_272 (.ZN (n_0_117), .A1 (hfn_ipo_n77), .A2 (n_0_155), .B1 (hfn_ipo_n75), .B2 (n_0_118));
OAI22_X1 i_0_271 (.ZN (n_0_116), .A1 (hfn_ipo_n67), .A2 (n_0_117), .B1 (hfn_ipo_n65), .B2 (n_0_137));
AOI22_X1 i_0_270 (.ZN (n_0_115), .A1 (hfn_ipo_n71), .A2 (n_0_126), .B1 (hfn_ipo_n69), .B2 (n_0_116));
OAI22_X1 i_0_269 (.ZN (n_0_114), .A1 (hfn_ipo_n79), .A2 (n_0_120), .B1 (hfn_ipo_n95), .B2 (n_0_115));
AND2_X1 i_0_268 (.ZN (n_284), .A1 (n_0_298), .A2 (n_0_114));
NOR2_X1 i_0_267 (.ZN (n_0_113), .A1 (n_0_380), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_266 (.ZN (n_0_112), .A1 (hfn_ipo_n77), .A2 (n_0_151), .B1 (hfn_ipo_n75), .B2 (n_0_113));
OAI22_X1 i_0_265 (.ZN (n_0_111), .A1 (hfn_ipo_n67), .A2 (n_0_112), .B1 (hfn_ipo_n65), .B2 (n_0_132));
AOI22_X1 i_0_264 (.ZN (n_0_110), .A1 (hfn_ipo_n69), .A2 (n_0_111), .B1 (hfn_ipo_n71), .B2 (n_0_121));
OAI22_X1 i_0_263 (.ZN (n_0_109), .A1 (hfn_ipo_n79), .A2 (n_0_115), .B1 (hfn_ipo_n94), .B2 (n_0_110));
AND2_X1 i_0_262 (.ZN (n_283), .A1 (n_0_298), .A2 (n_0_109));
NOR2_X1 i_0_261 (.ZN (n_0_108), .A1 (n_0_379), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_260 (.ZN (n_0_107), .A1 (hfn_ipo_n77), .A2 (n_0_147), .B1 (hfn_ipo_n75), .B2 (n_0_108));
OAI22_X1 i_0_259 (.ZN (n_0_106), .A1 (hfn_ipo_n67), .A2 (n_0_107), .B1 (hfn_ipo_n65), .B2 (n_0_127));
AOI22_X1 i_0_258 (.ZN (n_0_105), .A1 (hfn_ipo_n69), .A2 (n_0_106), .B1 (hfn_ipo_n71), .B2 (n_0_116));
OAI22_X1 i_0_257 (.ZN (n_0_104), .A1 (hfn_ipo_n94), .A2 (n_0_105), .B1 (hfn_ipo_n79), .B2 (n_0_110));
AND2_X1 i_0_256 (.ZN (n_282), .A1 (n_0_298), .A2 (n_0_104));
NOR2_X1 i_0_255 (.ZN (n_0_103), .A1 (n_0_378), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_254 (.ZN (n_0_102), .A1 (hfn_ipo_n75), .A2 (n_0_103), .B1 (hfn_ipo_n77), .B2 (n_0_143));
OAI22_X1 i_0_253 (.ZN (n_0_101), .A1 (hfn_ipo_n67), .A2 (n_0_102), .B1 (hfn_ipo_n65), .B2 (n_0_122));
AOI22_X1 i_0_252 (.ZN (n_0_100), .A1 (hfn_ipo_n69), .A2 (n_0_101), .B1 (hfn_ipo_n71), .B2 (n_0_111));
OAI22_X1 i_0_251 (.ZN (n_0_99), .A1 (hfn_ipo_n79), .A2 (n_0_105), .B1 (hfn_ipo_n94), .B2 (n_0_100));
AND2_X1 i_0_250 (.ZN (n_281), .A1 (n_0_298), .A2 (n_0_99));
NOR2_X1 i_0_249 (.ZN (n_0_98), .A1 (n_0_377), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_248 (.ZN (n_0_97), .A1 (hfn_ipo_n75), .A2 (n_0_98), .B1 (hfn_ipo_n77), .B2 (n_0_138));
OAI22_X1 i_0_247 (.ZN (n_0_96), .A1 (hfn_ipo_n65), .A2 (n_0_117), .B1 (hfn_ipo_n67), .B2 (n_0_97));
AOI22_X1 i_0_246 (.ZN (n_0_95), .A1 (hfn_ipo_n71), .A2 (n_0_106), .B1 (hfn_ipo_n69), .B2 (n_0_96));
OAI22_X1 i_0_245 (.ZN (n_0_94), .A1 (hfn_ipo_n79), .A2 (n_0_100), .B1 (hfn_ipo_n94), .B2 (n_0_95));
AND2_X1 i_0_244 (.ZN (n_280), .A1 (n_0_298), .A2 (n_0_94));
NOR2_X1 i_0_243 (.ZN (n_0_93), .A1 (n_0_376), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_242 (.ZN (n_0_92), .A1 (hfn_ipo_n75), .A2 (n_0_93), .B1 (hfn_ipo_n77), .B2 (n_0_133));
OAI22_X1 i_0_241 (.ZN (n_0_91), .A1 (hfn_ipo_n65), .A2 (n_0_112), .B1 (hfn_ipo_n67), .B2 (n_0_92));
AOI22_X1 i_0_240 (.ZN (n_0_90), .A1 (hfn_ipo_n71), .A2 (n_0_101), .B1 (hfn_ipo_n69), .B2 (n_0_91));
OAI22_X1 i_0_239 (.ZN (n_0_89), .A1 (hfn_ipo_n94), .A2 (n_0_90), .B1 (hfn_ipo_n79), .B2 (n_0_95));
AND2_X1 i_0_238 (.ZN (n_279), .A1 (n_0_298), .A2 (n_0_89));
NOR2_X1 i_0_237 (.ZN (n_0_88), .A1 (n_0_375), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_236 (.ZN (n_0_87), .A1 (hfn_ipo_n75), .A2 (n_0_88), .B1 (hfn_ipo_n77), .B2 (n_0_128));
OAI22_X1 i_0_235 (.ZN (n_0_86), .A1 (hfn_ipo_n65), .A2 (n_0_107), .B1 (hfn_ipo_n67), .B2 (n_0_87));
AOI22_X1 i_0_234 (.ZN (n_0_85), .A1 (hfn_ipo_n69), .A2 (n_0_86), .B1 (hfn_ipo_n71), .B2 (n_0_96));
OAI22_X1 i_0_233 (.ZN (n_0_84), .A1 (hfn_ipo_n79), .A2 (n_0_90), .B1 (hfn_ipo_n94), .B2 (n_0_85));
AND2_X1 i_0_232 (.ZN (n_278), .A1 (n_0_298), .A2 (n_0_84));
NOR2_X1 i_0_231 (.ZN (n_0_83), .A1 (n_0_374), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_230 (.ZN (n_0_82), .A1 (hfn_ipo_n75), .A2 (n_0_83), .B1 (hfn_ipo_n77), .B2 (n_0_123));
OAI22_X1 i_0_229 (.ZN (n_0_81), .A1 (hfn_ipo_n65), .A2 (n_0_102), .B1 (hfn_ipo_n67), .B2 (n_0_82));
AOI22_X1 i_0_228 (.ZN (n_0_80), .A1 (hfn_ipo_n69), .A2 (n_0_81), .B1 (hfn_ipo_n71), .B2 (n_0_91));
OAI22_X1 i_0_227 (.ZN (n_0_79), .A1 (hfn_ipo_n79), .A2 (n_0_85), .B1 (hfn_ipo_n94), .B2 (n_0_80));
AND2_X1 i_0_226 (.ZN (n_277), .A1 (n_0_298), .A2 (n_0_79));
NOR2_X1 i_0_225 (.ZN (n_0_78), .A1 (n_0_373), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_224 (.ZN (n_0_77), .A1 (hfn_ipo_n75), .A2 (n_0_78), .B1 (hfn_ipo_n77), .B2 (n_0_118));
OAI22_X1 i_0_223 (.ZN (n_0_76), .A1 (hfn_ipo_n67), .A2 (n_0_77), .B1 (hfn_ipo_n65), .B2 (n_0_97));
AOI22_X1 i_0_222 (.ZN (n_0_75), .A1 (hfn_ipo_n69), .A2 (n_0_76), .B1 (hfn_ipo_n71), .B2 (n_0_86));
OAI22_X1 i_0_221 (.ZN (n_0_74), .A1 (hfn_ipo_n94), .A2 (n_0_75), .B1 (hfn_ipo_n79), .B2 (n_0_80));
AND2_X1 i_0_220 (.ZN (n_276), .A1 (n_0_298), .A2 (n_0_74));
NOR2_X1 i_0_219 (.ZN (n_0_73), .A1 (n_0_372), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_218 (.ZN (n_0_72), .A1 (hfn_ipo_n75), .A2 (n_0_73), .B1 (hfn_ipo_n77), .B2 (n_0_113));
OAI22_X1 i_0_217 (.ZN (n_0_71), .A1 (hfn_ipo_n67), .A2 (n_0_72), .B1 (hfn_ipo_n65), .B2 (n_0_92));
AOI22_X1 i_0_216 (.ZN (n_0_70), .A1 (hfn_ipo_n71), .A2 (n_0_81), .B1 (hfn_ipo_n69), .B2 (n_0_71));
OAI22_X1 i_0_215 (.ZN (n_0_69), .A1 (hfn_ipo_n94), .A2 (n_0_70), .B1 (hfn_ipo_n79), .B2 (n_0_75));
AND2_X1 i_0_214 (.ZN (n_275), .A1 (n_0_298), .A2 (n_0_69));
NOR2_X1 i_0_213 (.ZN (n_0_68), .A1 (n_0_371), .A2 (hfn_ipo_n81));
AOI22_X1 i_0_212 (.ZN (n_0_67), .A1 (hfn_ipo_n75), .A2 (n_0_68), .B1 (hfn_ipo_n77), .B2 (n_0_108));
OAI22_X1 i_0_211 (.ZN (n_0_66), .A1 (hfn_ipo_n67), .A2 (n_0_67), .B1 (hfn_ipo_n65), .B2 (n_0_87));
AOI22_X1 i_0_210 (.ZN (n_0_65), .A1 (hfn_ipo_n69), .A2 (n_0_66), .B1 (hfn_ipo_n71), .B2 (n_0_76));
OAI22_X1 i_0_209 (.ZN (n_0_64), .A1 (hfn_ipo_n94), .A2 (n_0_65), .B1 (hfn_ipo_n79), .B2 (n_0_70));
AND2_X1 i_0_208 (.ZN (n_274), .A1 (n_0_298), .A2 (n_0_64));
AND2_X1 i_0_207 (.ZN (n_0_63), .A1 (n_357), .A2 (hfn_ipo_n83));
AOI22_X1 i_0_206 (.ZN (n_0_62), .A1 (hfn_ipo_n77), .A2 (n_0_103), .B1 (hfn_ipo_n75), .B2 (n_0_63));
OAI22_X1 i_0_205 (.ZN (n_0_61), .A1 (hfn_ipo_n65), .A2 (n_0_82), .B1 (hfn_ipo_n67), .B2 (n_0_62));
AOI22_X1 i_0_204 (.ZN (n_0_60), .A1 (hfn_ipo_n71), .A2 (n_0_71), .B1 (hfn_ipo_n69), .B2 (n_0_61));
OAI22_X1 i_0_203 (.ZN (n_0_59), .A1 (hfn_ipo_n79), .A2 (n_0_65), .B1 (hfn_ipo_n94), .B2 (n_0_60));
AND2_X1 i_0_202 (.ZN (n_273), .A1 (n_0_298), .A2 (n_0_59));
AND2_X1 i_0_201 (.ZN (n_0_58), .A1 (hfn_ipo_n77), .A2 (n_0_98));
NAND2_X1 i_0_200 (.ZN (n_0_57), .A1 (hfn_ipo_n65), .A2 (n_0_58));
OAI21_X1 i_0_199 (.ZN (n_0_56), .A (n_0_57), .B1 (hfn_ipo_n65), .B2 (n_0_77));
AOI22_X1 i_0_198 (.ZN (n_0_55), .A1 (hfn_ipo_n71), .A2 (n_0_66), .B1 (hfn_ipo_n69), .B2 (n_0_56));
OAI22_X1 i_0_197 (.ZN (n_0_54), .A1 (hfn_ipo_n79), .A2 (n_0_60), .B1 (hfn_ipo_n94), .B2 (n_0_55));
AND2_X1 i_0_196 (.ZN (n_272), .A1 (n_0_298), .A2 (n_0_54));
AND2_X1 i_0_195 (.ZN (n_0_53), .A1 (hfn_ipo_n77), .A2 (n_0_93));
NAND2_X1 i_0_194 (.ZN (n_0_52), .A1 (hfn_ipo_n65), .A2 (n_0_53));
OAI21_X1 i_0_193 (.ZN (n_0_51), .A (n_0_52), .B1 (hfn_ipo_n65), .B2 (n_0_72));
AOI22_X1 i_0_192 (.ZN (n_0_50), .A1 (hfn_ipo_n71), .A2 (n_0_61), .B1 (hfn_ipo_n69), .B2 (n_0_51));
OAI22_X1 i_0_191 (.ZN (n_0_49), .A1 (hfn_ipo_n79), .A2 (n_0_55), .B1 (hfn_ipo_n94), .B2 (n_0_50));
AND2_X1 i_0_190 (.ZN (n_271), .A1 (n_0_298), .A2 (n_0_49));
AND2_X1 i_0_189 (.ZN (n_0_48), .A1 (hfn_ipo_n77), .A2 (n_0_88));
NAND2_X1 i_0_188 (.ZN (n_0_47), .A1 (hfn_ipo_n65), .A2 (n_0_48));
OAI21_X1 i_0_187 (.ZN (n_0_46), .A (n_0_47), .B1 (hfn_ipo_n65), .B2 (n_0_67));
AOI22_X1 i_0_186 (.ZN (n_0_45), .A1 (hfn_ipo_n69), .A2 (n_0_46), .B1 (hfn_ipo_n71), .B2 (n_0_56));
OAI22_X1 i_0_185 (.ZN (n_0_44), .A1 (hfn_ipo_n79), .A2 (n_0_50), .B1 (hfn_ipo_n94), .B2 (n_0_45));
AND2_X1 i_0_184 (.ZN (n_270), .A1 (n_0_298), .A2 (n_0_44));
AND2_X1 i_0_183 (.ZN (n_0_43), .A1 (hfn_ipo_n77), .A2 (n_0_83));
NAND2_X1 i_0_182 (.ZN (n_0_42), .A1 (hfn_ipo_n65), .A2 (n_0_43));
OAI21_X1 i_0_181 (.ZN (n_0_41), .A (n_0_42), .B1 (hfn_ipo_n65), .B2 (n_0_62));
AOI22_X1 i_0_180 (.ZN (n_0_40), .A1 (hfn_ipo_n71), .A2 (n_0_51), .B1 (hfn_ipo_n69), .B2 (n_0_41));
OAI22_X1 i_0_179 (.ZN (n_0_39), .A1 (hfn_ipo_n79), .A2 (n_0_45), .B1 (hfn_ipo_n94), .B2 (n_0_40));
AND2_X1 i_0_178 (.ZN (n_269), .A1 (n_0_298), .A2 (n_0_39));
AND2_X1 i_0_177 (.ZN (n_0_38), .A1 (hfn_ipo_n77), .A2 (n_0_78));
AOI22_X1 i_0_176 (.ZN (n_0_37), .A1 (hfn_ipo_n65), .A2 (n_0_38), .B1 (hfn_ipo_n67), .B2 (n_0_58));
NAND2_X1 i_0_175 (.ZN (n_0_36), .A1 (hfn_ipo_n71), .A2 (n_0_46));
OAI21_X1 i_0_174 (.ZN (n_0_35), .A (n_0_36), .B1 (hfn_ipo_n71), .B2 (n_0_37));
NAND2_X1 i_0_173 (.ZN (n_0_34), .A1 (hfn_ipo_n79), .A2 (n_0_35));
OAI21_X1 i_0_172 (.ZN (n_0_33), .A (n_0_34), .B1 (hfn_ipo_n79), .B2 (n_0_40));
AND2_X1 i_0_171 (.ZN (n_268), .A1 (n_0_298), .A2 (n_0_33));
AND2_X1 i_0_170 (.ZN (n_0_32), .A1 (hfn_ipo_n77), .A2 (n_0_73));
AOI22_X1 i_0_169 (.ZN (n_0_31), .A1 (hfn_ipo_n65), .A2 (n_0_32), .B1 (hfn_ipo_n67), .B2 (n_0_53));
NAND2_X1 i_0_168 (.ZN (n_0_30), .A1 (hfn_ipo_n71), .A2 (n_0_41));
OAI21_X1 i_0_167 (.ZN (n_0_29), .A (n_0_30), .B1 (hfn_ipo_n71), .B2 (n_0_31));
AOI22_X1 i_0_166 (.ZN (n_0_28), .A1 (hfn_ipo_n94), .A2 (n_0_35), .B1 (hfn_ipo_n79), .B2 (n_0_29));
NOR2_X1 i_0_165 (.ZN (n_267), .A1 (drc_ipo_n96), .A2 (n_0_28));
AND2_X1 i_0_164 (.ZN (n_0_27), .A1 (hfn_ipo_n77), .A2 (n_0_68));
AOI22_X1 i_0_163 (.ZN (n_0_26), .A1 (hfn_ipo_n65), .A2 (n_0_27), .B1 (hfn_ipo_n67), .B2 (n_0_48));
OAI22_X1 i_0_162 (.ZN (n_0_25), .A1 (hfn_ipo_n71), .A2 (n_0_26), .B1 (hfn_ipo_n69), .B2 (n_0_37));
AOI22_X1 i_0_161 (.ZN (n_0_24), .A1 (hfn_ipo_n94), .A2 (n_0_29), .B1 (hfn_ipo_n79), .B2 (n_0_25));
NOR2_X1 i_0_160 (.ZN (n_266), .A1 (drc_ipo_n96), .A2 (n_0_24));
AND2_X1 i_0_159 (.ZN (n_0_23), .A1 (hfn_ipo_n77), .A2 (n_0_63));
AOI22_X1 i_0_158 (.ZN (n_0_22), .A1 (hfn_ipo_n67), .A2 (n_0_43), .B1 (hfn_ipo_n65), .B2 (n_0_23));
OAI22_X1 i_0_157 (.ZN (n_0_21), .A1 (hfn_ipo_n69), .A2 (n_0_31), .B1 (hfn_ipo_n71), .B2 (n_0_22));
AOI22_X1 i_0_156 (.ZN (n_0_20), .A1 (hfn_ipo_n94), .A2 (n_0_25), .B1 (hfn_ipo_n79), .B2 (n_0_21));
NOR2_X1 i_0_155 (.ZN (n_265), .A1 (drc_ipo_n96), .A2 (n_0_20));
AND2_X1 i_0_154 (.ZN (n_0_19), .A1 (hfn_ipo_n67), .A2 (n_0_38));
NAND2_X1 i_0_153 (.ZN (n_0_18), .A1 (hfn_ipo_n69), .A2 (n_0_19));
OAI21_X1 i_0_152 (.ZN (n_0_17), .A (n_0_18), .B1 (hfn_ipo_n69), .B2 (n_0_26));
AOI22_X1 i_0_151 (.ZN (n_0_16), .A1 (hfn_ipo_n94), .A2 (n_0_21), .B1 (hfn_ipo_n79), .B2 (n_0_17));
NOR2_X1 i_0_150 (.ZN (n_264), .A1 (drc_ipo_n96), .A2 (n_0_16));
AND2_X1 i_0_149 (.ZN (n_0_15), .A1 (hfn_ipo_n67), .A2 (n_0_32));
NAND2_X1 i_0_148 (.ZN (n_0_14), .A1 (hfn_ipo_n69), .A2 (n_0_15));
OAI21_X1 i_0_147 (.ZN (n_0_13), .A (n_0_14), .B1 (hfn_ipo_n69), .B2 (n_0_22));
AOI22_X1 i_0_146 (.ZN (n_0_12), .A1 (hfn_ipo_n94), .A2 (n_0_17), .B1 (hfn_ipo_n79), .B2 (n_0_13));
NOR2_X1 i_0_145 (.ZN (n_263), .A1 (drc_ipo_n96), .A2 (n_0_12));
NAND2_X1 i_0_144 (.ZN (n_0_11), .A1 (hfn_ipo_n94), .A2 (n_0_13));
AND2_X1 i_0_143 (.ZN (n_0_10), .A1 (hfn_ipo_n67), .A2 (n_0_27));
AOI22_X1 i_0_142 (.ZN (n_0_9), .A1 (hfn_ipo_n69), .A2 (n_0_10), .B1 (hfn_ipo_n71), .B2 (n_0_19));
OR2_X1 i_0_141 (.ZN (n_0_8), .A1 (hfn_ipo_n94), .A2 (n_0_9));
AOI21_X1 i_0_140 (.ZN (n_262), .A (drc_ipo_n96), .B1 (n_0_11), .B2 (n_0_8));
AND2_X1 i_0_139 (.ZN (n_0_7), .A1 (hfn_ipo_n67), .A2 (n_0_23));
AOI22_X1 i_0_138 (.ZN (n_0_6), .A1 (hfn_ipo_n71), .A2 (n_0_15), .B1 (hfn_ipo_n69), .B2 (n_0_7));
OAI22_X1 i_0_137 (.ZN (n_0_5), .A1 (hfn_ipo_n79), .A2 (n_0_9), .B1 (hfn_ipo_n94), .B2 (n_0_6));
AND2_X1 i_0_136 (.ZN (n_261), .A1 (n_0_298), .A2 (n_0_5));
NAND2_X1 i_0_135 (.ZN (n_0_4), .A1 (hfn_ipo_n71), .A2 (n_0_10));
AOI221_X1 i_0_134 (.ZN (n_260), .A (drc_ipo_n96), .B1 (hfn_ipo_n94), .B2 (n_0_6), .C1 (hfn_ipo_n79), .C2 (n_0_4));
NAND2_X1 i_0_133 (.ZN (n_0_3), .A1 (hfn_ipo_n71), .A2 (n_0_7));
AOI221_X1 i_0_132 (.ZN (n_259), .A (drc_ipo_n96), .B1 (hfn_ipo_n94), .B2 (n_0_4), .C1 (hfn_ipo_n79), .C2 (n_0_3));
NOR3_X1 i_0_131 (.ZN (n_258), .A1 (hfn_ipo_n79), .A2 (n_0_3), .A3 (drc_ipo_n96));
AND2_X1 i_0_130 (.ZN (n_257), .A1 (n_0_442), .A2 (\acc_out[63] ));
AND2_X1 i_0_129 (.ZN (n_256), .A1 (n_0_442), .A2 (\acc_out[62] ));
AND2_X1 i_0_128 (.ZN (n_255), .A1 (n_0_442), .A2 (\acc_out[61] ));
AND2_X1 i_0_127 (.ZN (n_254), .A1 (n_0_442), .A2 (\acc_out[60] ));
AND2_X1 i_0_126 (.ZN (n_253), .A1 (n_0_442), .A2 (\acc_out[59] ));
AND2_X1 i_0_125 (.ZN (n_252), .A1 (n_0_442), .A2 (\acc_out[58] ));
AND2_X1 i_0_124 (.ZN (n_251), .A1 (n_0_442), .A2 (\acc_out[57] ));
AND2_X1 i_0_123 (.ZN (n_250), .A1 (n_0_442), .A2 (\acc_out[56] ));
AND2_X1 i_0_122 (.ZN (n_249), .A1 (n_0_442), .A2 (\acc_out[55] ));
AND2_X1 i_0_121 (.ZN (n_248), .A1 (n_0_442), .A2 (\acc_out[54] ));
AND2_X1 i_0_120 (.ZN (n_247), .A1 (n_0_442), .A2 (\acc_out[53] ));
AND2_X1 i_0_119 (.ZN (n_246), .A1 (n_0_442), .A2 (\acc_out[52] ));
AND2_X1 i_0_118 (.ZN (n_245), .A1 (n_0_442), .A2 (\acc_out[51] ));
AND2_X1 i_0_117 (.ZN (n_244), .A1 (n_0_442), .A2 (\acc_out[50] ));
AND2_X1 i_0_116 (.ZN (n_243), .A1 (hfn_ipo_n91), .A2 (\acc_out[49] ));
AND2_X1 i_0_115 (.ZN (n_242), .A1 (hfn_ipo_n91), .A2 (\acc_out[48] ));
AND2_X1 i_0_114 (.ZN (n_241), .A1 (hfn_ipo_n91), .A2 (\acc_out[47] ));
AND2_X1 i_0_113 (.ZN (n_240), .A1 (hfn_ipo_n91), .A2 (\acc_out[46] ));
AND2_X1 i_0_112 (.ZN (n_239), .A1 (hfn_ipo_n91), .A2 (\acc_out[45] ));
AND2_X1 i_0_111 (.ZN (n_238), .A1 (hfn_ipo_n91), .A2 (\acc_out[44] ));
AND2_X1 i_0_110 (.ZN (n_237), .A1 (hfn_ipo_n91), .A2 (\acc_out[43] ));
AND2_X1 i_0_109 (.ZN (n_236), .A1 (hfn_ipo_n91), .A2 (\acc_out[42] ));
AND2_X1 i_0_108 (.ZN (n_235), .A1 (hfn_ipo_n91), .A2 (\acc_out[41] ));
AND2_X1 i_0_107 (.ZN (n_234), .A1 (hfn_ipo_n91), .A2 (\acc_out[40] ));
AND2_X1 i_0_106 (.ZN (n_233), .A1 (hfn_ipo_n91), .A2 (\acc_out[39] ));
AND2_X1 i_0_105 (.ZN (n_232), .A1 (hfn_ipo_n91), .A2 (\acc_out[38] ));
AND2_X1 i_0_104 (.ZN (n_231), .A1 (hfn_ipo_n91), .A2 (\acc_out[37] ));
AND2_X1 i_0_103 (.ZN (n_230), .A1 (hfn_ipo_n91), .A2 (\acc_out[36] ));
AND2_X1 i_0_102 (.ZN (n_229), .A1 (hfn_ipo_n91), .A2 (\acc_out[35] ));
AND2_X1 i_0_101 (.ZN (n_228), .A1 (hfn_ipo_n91), .A2 (\acc_out[34] ));
AND2_X1 i_0_100 (.ZN (n_227), .A1 (hfn_ipo_n91), .A2 (\acc_out[33] ));
AND2_X1 i_0_99 (.ZN (n_226), .A1 (hfn_ipo_n91), .A2 (\acc_out[32] ));
AND2_X1 i_0_98 (.ZN (n_225), .A1 (hfn_ipo_n91), .A2 (\acc_out[31] ));
AND2_X1 i_0_97 (.ZN (n_224), .A1 (hfn_ipo_n91), .A2 (\acc_out[30] ));
AND2_X1 i_0_96 (.ZN (n_223), .A1 (hfn_ipo_n91), .A2 (\acc_out[29] ));
AND2_X1 i_0_95 (.ZN (n_222), .A1 (hfn_ipo_n91), .A2 (\acc_out[28] ));
AND2_X1 i_0_94 (.ZN (n_221), .A1 (hfn_ipo_n91), .A2 (\acc_out[27] ));
AND2_X1 i_0_93 (.ZN (n_220), .A1 (hfn_ipo_n91), .A2 (\acc_out[26] ));
AND2_X1 i_0_92 (.ZN (n_219), .A1 (hfn_ipo_n91), .A2 (\acc_out[25] ));
AND2_X1 i_0_91 (.ZN (n_218), .A1 (hfn_ipo_n91), .A2 (\acc_out[24] ));
AND2_X1 i_0_90 (.ZN (n_217), .A1 (hfn_ipo_n90), .A2 (\acc_out[23] ));
AND2_X1 i_0_89 (.ZN (n_216), .A1 (hfn_ipo_n90), .A2 (\acc_out[22] ));
AND2_X1 i_0_88 (.ZN (n_215), .A1 (hfn_ipo_n90), .A2 (\acc_out[21] ));
AND2_X1 i_0_87 (.ZN (n_214), .A1 (hfn_ipo_n90), .A2 (\acc_out[20] ));
AND2_X1 i_0_86 (.ZN (n_213), .A1 (hfn_ipo_n90), .A2 (\acc_out[19] ));
AND2_X1 i_0_85 (.ZN (n_212), .A1 (hfn_ipo_n90), .A2 (\acc_out[18] ));
AND2_X1 i_0_84 (.ZN (n_211), .A1 (hfn_ipo_n90), .A2 (\acc_out[17] ));
AND2_X1 i_0_83 (.ZN (n_210), .A1 (hfn_ipo_n90), .A2 (\acc_out[16] ));
AND2_X1 i_0_82 (.ZN (n_209), .A1 (hfn_ipo_n90), .A2 (\acc_out[15] ));
AND2_X1 i_0_81 (.ZN (n_208), .A1 (hfn_ipo_n90), .A2 (\acc_out[14] ));
AND2_X1 i_0_80 (.ZN (n_207), .A1 (hfn_ipo_n90), .A2 (\acc_out[13] ));
AND2_X1 i_0_79 (.ZN (n_206), .A1 (hfn_ipo_n90), .A2 (\acc_out[12] ));
AND2_X1 i_0_78 (.ZN (n_205), .A1 (hfn_ipo_n90), .A2 (\acc_out[11] ));
AND2_X1 i_0_77 (.ZN (n_204), .A1 (hfn_ipo_n90), .A2 (\acc_out[10] ));
AND2_X1 i_0_76 (.ZN (n_203), .A1 (hfn_ipo_n90), .A2 (\acc_out[9] ));
AND2_X1 i_0_75 (.ZN (n_202), .A1 (hfn_ipo_n90), .A2 (\acc_out[8] ));
AND2_X1 i_0_74 (.ZN (n_201), .A1 (hfn_ipo_n90), .A2 (\acc_out[7] ));
AND2_X1 i_0_73 (.ZN (n_200), .A1 (hfn_ipo_n90), .A2 (\acc_out[6] ));
AND2_X1 i_0_72 (.ZN (n_199), .A1 (hfn_ipo_n90), .A2 (\acc_out[5] ));
AND2_X1 i_0_71 (.ZN (n_198), .A1 (hfn_ipo_n90), .A2 (\acc_out[4] ));
AND2_X1 i_0_70 (.ZN (n_197), .A1 (hfn_ipo_n90), .A2 (\acc_out[3] ));
AND2_X1 i_0_69 (.ZN (n_196), .A1 (hfn_ipo_n90), .A2 (\acc_out[2] ));
AND2_X1 i_0_68 (.ZN (n_195), .A1 (hfn_ipo_n90), .A2 (\acc_out[1] ));
AND2_X1 i_0_67 (.ZN (n_194), .A1 (hfn_ipo_n90), .A2 (\acc_out[0] ));
AND2_X1 i_0_66 (.ZN (n_193), .A1 (n_126), .A2 (hfn_ipo_n73));
AND2_X1 i_0_65 (.ZN (n_192), .A1 (n_125), .A2 (hfn_ipo_n73));
AND2_X1 i_0_64 (.ZN (n_191), .A1 (n_124), .A2 (hfn_ipo_n73));
AND2_X1 i_0_63 (.ZN (n_190), .A1 (n_123), .A2 (hfn_ipo_n73));
AND2_X1 i_0_62 (.ZN (n_189), .A1 (n_122), .A2 (hfn_ipo_n73));
AND2_X1 i_0_61 (.ZN (n_188), .A1 (n_121), .A2 (hfn_ipo_n73));
AND2_X1 i_0_60 (.ZN (n_187), .A1 (n_120), .A2 (hfn_ipo_n73));
AND2_X1 i_0_59 (.ZN (n_186), .A1 (n_119), .A2 (hfn_ipo_n73));
AND2_X1 i_0_58 (.ZN (n_185), .A1 (n_118), .A2 (hfn_ipo_n73));
AND2_X1 i_0_57 (.ZN (n_184), .A1 (n_117), .A2 (hfn_ipo_n73));
AND2_X1 i_0_56 (.ZN (n_183), .A1 (n_116), .A2 (hfn_ipo_n73));
AND2_X1 i_0_55 (.ZN (n_182), .A1 (n_115), .A2 (hfn_ipo_n73));
AND2_X1 i_0_54 (.ZN (n_181), .A1 (n_114), .A2 (hfn_ipo_n73));
AND2_X1 i_0_53 (.ZN (n_180), .A1 (n_113), .A2 (hfn_ipo_n73));
AND2_X1 i_0_52 (.ZN (n_179), .A1 (n_112), .A2 (hfn_ipo_n73));
AND2_X1 i_0_51 (.ZN (n_178), .A1 (n_111), .A2 (hfn_ipo_n74));
AND2_X1 i_0_50 (.ZN (n_177), .A1 (n_110), .A2 (hfn_ipo_n74));
AND2_X1 i_0_49 (.ZN (n_176), .A1 (n_109), .A2 (hfn_ipo_n74));
AND2_X1 i_0_48 (.ZN (n_175), .A1 (n_108), .A2 (hfn_ipo_n74));
AND2_X1 i_0_47 (.ZN (n_174), .A1 (n_107), .A2 (hfn_ipo_n74));
AND2_X1 i_0_46 (.ZN (n_173), .A1 (n_106), .A2 (hfn_ipo_n74));
AND2_X1 i_0_45 (.ZN (n_172), .A1 (n_105), .A2 (hfn_ipo_n74));
AND2_X1 i_0_44 (.ZN (n_171), .A1 (n_104), .A2 (hfn_ipo_n74));
AND2_X1 i_0_43 (.ZN (n_170), .A1 (n_103), .A2 (hfn_ipo_n74));
AND2_X1 i_0_42 (.ZN (n_169), .A1 (n_102), .A2 (hfn_ipo_n74));
AND2_X1 i_0_41 (.ZN (n_168), .A1 (n_101), .A2 (hfn_ipo_n74));
AND2_X1 i_0_40 (.ZN (n_167), .A1 (n_100), .A2 (hfn_ipo_n74));
AND2_X1 i_0_39 (.ZN (n_166), .A1 (n_99), .A2 (hfn_ipo_n74));
AND2_X1 i_0_38 (.ZN (n_165), .A1 (n_98), .A2 (hfn_ipo_n74));
AND2_X1 i_0_37 (.ZN (n_164), .A1 (n_97), .A2 (hfn_ipo_n74));
AND2_X1 i_0_36 (.ZN (n_163), .A1 (n_96), .A2 (hfn_ipo_n74));
AND2_X1 i_0_35 (.ZN (n_162), .A1 (n_95), .A2 (hfn_ipo_n74));
AND2_X1 i_0_34 (.ZN (n_161), .A1 (n_94), .A2 (hfn_ipo_n74));
AND2_X1 i_0_33 (.ZN (n_160), .A1 (n_93), .A2 (hfn_ipo_n74));
AND2_X1 i_0_32 (.ZN (n_159), .A1 (n_92), .A2 (hfn_ipo_n74));
AND2_X1 i_0_31 (.ZN (n_158), .A1 (n_91), .A2 (hfn_ipo_n74));
AND2_X1 i_0_30 (.ZN (n_157), .A1 (n_90), .A2 (hfn_ipo_n74));
AND2_X1 i_0_29 (.ZN (n_156), .A1 (n_89), .A2 (hfn_ipo_n74));
AND2_X1 i_0_28 (.ZN (n_155), .A1 (n_88), .A2 (hfn_ipo_n74));
AND2_X1 i_0_27 (.ZN (n_154), .A1 (n_87), .A2 (hfn_ipo_n74));
AND2_X1 i_0_26 (.ZN (n_153), .A1 (n_86), .A2 (hfn_ipo_n73));
AND2_X1 i_0_25 (.ZN (n_152), .A1 (n_85), .A2 (hfn_ipo_n73));
AND2_X1 i_0_24 (.ZN (n_151), .A1 (n_84), .A2 (hfn_ipo_n73));
AND2_X1 i_0_23 (.ZN (n_150), .A1 (n_83), .A2 (hfn_ipo_n73));
AND2_X1 i_0_22 (.ZN (n_149), .A1 (n_82), .A2 (hfn_ipo_n73));
AND2_X1 i_0_21 (.ZN (n_148), .A1 (n_81), .A2 (hfn_ipo_n73));
AND2_X1 i_0_20 (.ZN (n_147), .A1 (n_80), .A2 (hfn_ipo_n73));
AND2_X1 i_0_19 (.ZN (n_146), .A1 (n_79), .A2 (hfn_ipo_n73));
AND2_X1 i_0_18 (.ZN (n_145), .A1 (n_78), .A2 (hfn_ipo_n73));
AND2_X1 i_0_17 (.ZN (n_144), .A1 (n_77), .A2 (hfn_ipo_n73));
AND2_X1 i_0_16 (.ZN (n_143), .A1 (n_76), .A2 (hfn_ipo_n73));
AND2_X1 i_0_15 (.ZN (n_142), .A1 (n_75), .A2 (hfn_ipo_n73));
AND2_X1 i_0_14 (.ZN (n_141), .A1 (n_74), .A2 (hfn_ipo_n73));
AND2_X1 i_0_13 (.ZN (n_140), .A1 (n_73), .A2 (hfn_ipo_n73));
AND2_X1 i_0_12 (.ZN (n_139), .A1 (n_72), .A2 (hfn_ipo_n73));
AND2_X1 i_0_11 (.ZN (n_138), .A1 (n_71), .A2 (hfn_ipo_n73));
AND2_X1 i_0_10 (.ZN (n_137), .A1 (n_70), .A2 (hfn_ipo_n73));
AND2_X1 i_0_9 (.ZN (n_136), .A1 (n_69), .A2 (hfn_ipo_n73));
AND2_X1 i_0_8 (.ZN (n_135), .A1 (n_68), .A2 (hfn_ipo_n73));
AND2_X1 i_0_7 (.ZN (n_134), .A1 (n_67), .A2 (hfn_ipo_n73));
AND2_X1 i_0_6 (.ZN (n_133), .A1 (n_66), .A2 (hfn_ipo_n73));
AND2_X1 i_0_5 (.ZN (n_132), .A1 (n_65), .A2 (hfn_ipo_n73));
AND2_X1 i_0_4 (.ZN (n_131), .A1 (n_64), .A2 (hfn_ipo_n73));
AND2_X1 i_0_3 (.ZN (n_130), .A1 (n_63), .A2 (hfn_ipo_n73));
HA_X1 i_0_2 (.CO (n_0_2), .S (n_129), .A (hfn_ipo_n75), .B (n_0_1));
HA_X1 i_0_1 (.CO (n_0_1), .S (n_128), .A (hfn_ipo_n65), .B (n_0_0));
HA_X1 i_0_0 (.CO (n_0_0), .S (n_127), .A (hfn_ipo_n69), .B (hfn_ipo_n79));
datapath__0_10 i_13 (.acc_out1 ({n_126, n_125, n_124, n_123, n_122, n_121, n_120, 
    n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, 
    n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63}), .acc_out ({n_257, n_256, n_255, 
    n_254, n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, 
    n_243, n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, 
    n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, 
    n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, 
    n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, 
    n_199, n_198, n_197, n_196, n_195, n_194}), .p_0 ({n_321, n_320, n_319, n_318, 
    n_317, n_316, n_315, n_314, n_313, n_312, n_311, n_310, n_309, n_308, n_307, 
    n_306, n_305, n_304, n_303, n_302, n_301, n_300, n_299, n_298, n_297, n_296, 
    n_295, n_294, n_293, n_292, n_291, n_290, n_289, n_288, n_287, n_286, n_285, 
    n_284, n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, 
    n_273, n_272, n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, 
    n_262, n_261, n_260, n_259, n_258}));
datapath__0_5 i_8 (.p_0 ({n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, uc_1}), .in2 ({in2[31], in2[30], 
    in2[29], in2[28], in2[27], in2[26], in2[25], in2[24], in2[23], in2[22], in2[21], 
    in2[20], in2[19], in2[18], in2[17], in2[16], in2[15], in2[14], in2[13], in2[12], 
    in2[11], in2[10], in2[9], in2[8], in2[7], in2[6], in2[5], in2[4], in2[3], in2[2], 
    in2[1], in2[0]}));
datapath i_2 (.p_0 ({n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, 
    n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, 
    n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, uc_0}), .in1 ({in1[31], in1[30], in1[29], 
    in1[28], in1[27], in1[26], in1[25], in1[24], in1[23], in1[22], in1[21], in1[20], 
    in1[19], in1[18], in1[17], in1[16], in1[15], in1[14], in1[13], in1[12], in1[11], 
    in1[10], in1[9], in1[8], in1[7], in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], 
    in1[0]}));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n105), .D (n_130));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n105), .D (n_131));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n105), .D (n_132));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n105), .D (n_133));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n105), .D (n_134));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n105), .D (n_135));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n105), .D (n_136));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n105), .D (n_137));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n105), .D (n_138));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n105), .D (n_139));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n105), .D (n_140));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n105), .D (n_141));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n105), .D (n_142));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n105), .D (n_143));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n105), .D (n_144));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n105), .D (n_145));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n105), .D (n_146));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n105), .D (n_147));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n105), .D (n_148));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n105), .D (n_149));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n105), .D (n_150));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n105), .D (n_151));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n105), .D (n_152));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n105), .D (n_153));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n105), .D (n_154));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n105), .D (n_155));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n105), .D (n_156));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n105), .D (n_157));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n105), .D (n_158));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n105), .D (n_159));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n105), .D (n_160));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n105), .D (n_161));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n105), .D (n_162));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n105), .D (n_163));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n105), .D (n_164));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n105), .D (n_165));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n105), .D (n_166));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n105), .D (n_167));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n105), .D (n_168));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n105), .D (n_169));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n105), .D (n_170));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (CTS_n105), .D (n_171));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (CTS_n105), .D (n_172));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (CTS_n105), .D (n_173));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (CTS_n105), .D (n_174));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (CTS_n105), .D (n_175));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (CTS_n105), .D (n_176));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (CTS_n105), .D (n_177));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (CTS_n105), .D (n_178));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (CTS_n105), .D (n_179));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (CTS_n105), .D (n_180));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (CTS_n105), .D (n_181));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (CTS_n105), .D (n_182));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (CTS_n105), .D (n_183));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (CTS_n105), .D (n_184));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (CTS_n105), .D (n_185));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (CTS_n105), .D (n_186));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (CTS_n105), .D (n_187));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (CTS_n105), .D (n_188));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (CTS_n105), .D (n_189));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (CTS_n105), .D (n_190));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (CTS_n105), .D (n_191));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (CTS_n105), .D (n_192));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (CTS_n105), .D (n_193));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n106), .CK (clk_CTSPP_236), .E (n_354), .SE (1'b0 ));
BUF_X2 hfn_ipo_c72 (.Z (hfn_ipo_n72), .A (n_0_330));
BUF_X4 hfn_ipo_c73 (.Z (hfn_ipo_n73), .A (n_0_363));
BUF_X2 hfn_ipo_c71 (.Z (hfn_ipo_n71), .A (n_0_330));
CLKBUF_X1 hfn_ipo_c74 (.Z (hfn_ipo_n74), .A (n_0_363));
BUF_X2 hfn_ipo_c76 (.Z (hfn_ipo_n76), .A (n_0_365));
CLKBUF_X1 hfn_ipo_c77 (.Z (hfn_ipo_n77), .A (n_0_366));
BUF_X2 hfn_ipo_c75 (.Z (hfn_ipo_n75), .A (n_0_365));
CLKBUF_X1 hfn_ipo_c78 (.Z (hfn_ipo_n78), .A (n_0_366));
BUF_X4 hfn_ipo_c79 (.Z (hfn_ipo_n79), .A (n_0_367));
BUF_X2 hfn_ipo_c80 (.Z (hfn_ipo_n80), .A (n_0_367));
CLKBUF_X2 hfn_ipo_c82 (.Z (hfn_ipo_n82), .A (n_0_368));
CLKBUF_X1 hfn_ipo_c83 (.Z (hfn_ipo_n83), .A (n_0_369));
CLKBUF_X2 hfn_ipo_c81 (.Z (hfn_ipo_n81), .A (n_0_368));
CLKBUF_X3 CTS_L3_c106 (.Z (CTS_n105), .A (CTS_n106));
BUF_X2 hfn_ipo_c94 (.Z (hfn_ipo_n94), .A (n_355));
BUF_X2 hfn_ipo_c95 (.Z (hfn_ipo_n95), .A (n_355));
CLKBUF_X2 hfn_ipo_c86 (.Z (hfn_ipo_n86), .A (n_0_436));
CLKBUF_X2 hfn_ipo_c87 (.Z (hfn_ipo_n87), .A (n_0_438));
CLKBUF_X2 hfn_ipo_c85 (.Z (hfn_ipo_n85), .A (n_0_436));
CLKBUF_X2 hfn_ipo_c88 (.Z (hfn_ipo_n88), .A (n_0_438));
BUF_X4 hfn_ipo_c89 (.Z (hfn_ipo_n89), .A (n_0_442));
CLKBUF_X1 hfn_ipo_c90 (.Z (hfn_ipo_n90), .A (n_0_442));
BUF_X2 hfn_ipo_c91 (.Z (hfn_ipo_n91), .A (n_0_442));
CLKBUF_X1 hfn_ipo_c92 (.Z (hfn_ipo_n92), .A (n_0_442));
BUF_X2 hfn_ipo_c65 (.Z (hfn_ipo_n65), .A (n_0_327));
BUF_X2 hfn_ipo_c66 (.Z (hfn_ipo_n66), .A (n_0_327));
CLKBUF_X2 hfn_ipo_c67 (.Z (hfn_ipo_n67), .A (n_0_328));
CLKBUF_X2 hfn_ipo_c68 (.Z (hfn_ipo_n68), .A (n_0_328));
BUF_X4 hfn_ipo_c69 (.Z (hfn_ipo_n69), .A (n_0_329));
BUF_X4 drc_ipo_c96 (.Z (drc_ipo_n96), .A (n_0_299));
BUF_X2 hfn_ipo_c70 (.Z (hfn_ipo_n70), .A (n_0_329));
CLKBUF_X1 CLOCK_slh__c236 (.Z (n_322), .A (CLOCK_slh__n1277));
CLKBUF_X3 CTS_L2_c233 (.Z (clk_CTSPP_233), .A (clk_CTSPP_236));

endmodule //sequential_multiplier

module Register (clk_CTSPP_119, clk_CTSPP_120, clk_CTSPP_122, clk_CTSPP_125, in, 
    clk, out);

output [31:0] out;
output clk_CTSPP_119;
output clk_CTSPP_120;
input clk;
input [31:0] in;
input clk_CTSPP_122;
input clk_CTSPP_125;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk_CTSPP_120), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk_CTSPP_120), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk_CTSPP_119), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk_CTSPP_119), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk_CTSPP_119), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk_CTSPP_119), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk_CTSPP_119), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk_CTSPP_122), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk_CTSPP_122), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk_CTSPP_122), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk_CTSPP_122), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk_CTSPP_119), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk_CTSPP_119), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk_CTSPP_119), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk_CTSPP_119), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk_CTSPP_119), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk_CTSPP_119), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk_CTSPP_119), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk_CTSPP_119), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk_CTSPP_119), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk_CTSPP_119), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk_CTSPP_119), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk_CTSPP_119), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk_CTSPP_119), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk_CTSPP_120), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk_CTSPP_119), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk_CTSPP_119), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk_CTSPP_119), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk_CTSPP_120), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk_CTSPP_120), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk_CTSPP_120), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk_CTSPP_120), .D (in[31]));
CLKBUF_X2 CTS_L2_c50 (.Z (clk_CTSPP_120), .A (clk_CTSPP_125));
CLKBUF_X2 CTS_L2_c48 (.Z (clk_CTSPP_119), .A (clk_CTSPP_125));

endmodule //Register

module Register__0_13 (clk_CTSPP_192, clk_CTSPP_191, clk_CTSPP_193, clk_CTSPP_195, 
    clk_CTSPP_196, clk_CTSPP_198, in, clk, out);

output [31:0] out;
output clk_CTSPP_192;
input clk;
input [31:0] in;
input clk_CTSPP_191;
input clk_CTSPP_193;
input clk_CTSPP_195;
input clk_CTSPP_196;
input clk_CTSPP_198;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk_CTSPP_195), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk_CTSPP_195), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk_CTSPP_195), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk_CTSPP_195), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk_CTSPP_195), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk_CTSPP_191), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk_CTSPP_191), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk_CTSPP_195), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk_CTSPP_195), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk_CTSPP_196), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk_CTSPP_195), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk_CTSPP_193), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk_CTSPP_193), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk_CTSPP_192), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk_CTSPP_193), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk_CTSPP_193), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk_CTSPP_193), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk_CTSPP_193), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk_CTSPP_193), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk_CTSPP_193), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk_CTSPP_193), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk_CTSPP_193), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk_CTSPP_193), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk_CTSPP_193), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk_CTSPP_193), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk_CTSPP_193), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk_CTSPP_193), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk_CTSPP_193), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk_CTSPP_192), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk_CTSPP_192), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk_CTSPP_192), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk_CTSPP_193), .D (in[31]));
CLKBUF_X2 CTS_L2_c18 (.Z (clk_CTSPP_192), .A (clk_CTSPP_198));

endmodule //Register__0_13

module SequentialMultiplierIntegerated (in1, in2, clk, rst, out);

output [63:0] out;
input clk;
input [31:0] in1;
input [31:0] in2;
input rst;
wire CLOCK_slh_n869;
wire CLOCK_slh_n944;
wire CLOCK_slh_n939;
wire CLOCK_slh_n949;
wire CLOCK_slh_n934;
wire CLOCK_slh_n929;
wire CLOCK_slh_n879;
wire CLOCK_slh_n904;
wire CLOCK_slh_n874;
wire CLOCK_slh_n854;
wire CLOCK_slh_n899;
wire CLOCK_slh_n894;
wire CLOCK_slh_n849;
wire CLOCK_slh_n839;
wire CLOCK_slh_n859;
wire CLOCK_slh_n819;
wire CLOCK_slh_n834;
wire CLOCK_slh_n919;
wire CLOCK_slh_n924;
wire CLOCK_slh_n829;
wire CLOCK_slh_n814;
wire CLOCK_slh_n954;
wire CLOCK_slh_n699;
wire CLOCK_slh_n704;
wire CLOCK_slh_n824;
wire CLOCK_slh_n844;
wire CLOCK_slh_n914;
wire CLOCK_slh_n909;
wire CLOCK_slh_n804;
wire CLOCK_slh_n754;
wire CLOCK_slh_n799;
wire CLOCK_slh_n889;
wire CLOCK_slh_n794;
wire CLOCK_slh_n789;
wire CLOCK_slh_n784;
wire CLOCK_slh_n779;
wire CLOCK_slh_n774;
wire CLOCK_slh_n769;
wire CLOCK_slh_n764;
wire CLOCK_slh_n759;
wire CLOCK_slh_n744;
wire CLOCK_slh_n749;
wire CLOCK_slh_n739;
wire CLOCK_slh_n734;
wire CLOCK_slh_n729;
wire CLOCK_slh_n719;
wire CLOCK_slh_n724;
wire CLOCK_slh_n709;
wire CLOCK_slh_n714;
wire CLOCK_slh_n809;
wire CLOCK_slh_n884;
wire CLOCK_slh_n864;
wire \operand1[31] ;
wire \operand1[30] ;
wire \operand1[29] ;
wire \operand1[28] ;
wire \operand1[27] ;
wire \operand1[26] ;
wire \operand1[25] ;
wire \operand1[24] ;
wire \operand1[23] ;
wire \operand1[22] ;
wire \operand1[21] ;
wire \operand1[20] ;
wire \operand1[19] ;
wire \operand1[18] ;
wire \operand1[17] ;
wire \operand1[16] ;
wire \operand1[15] ;
wire \operand1[14] ;
wire \operand1[13] ;
wire \operand1[12] ;
wire \operand1[11] ;
wire \operand1[10] ;
wire \operand1[9] ;
wire \operand1[8] ;
wire \operand1[7] ;
wire \operand1[6] ;
wire \operand1[5] ;
wire \operand1[4] ;
wire \operand1[3] ;
wire \operand1[2] ;
wire \operand1[1] ;
wire \operand1[0] ;
wire \operand2[31] ;
wire \operand2[30] ;
wire \operand2[29] ;
wire \operand2[28] ;
wire \operand2[27] ;
wire \operand2[26] ;
wire \operand2[25] ;
wire \operand2[24] ;
wire \operand2[23] ;
wire \operand2[22] ;
wire \operand2[21] ;
wire \operand2[20] ;
wire \operand2[19] ;
wire \operand2[18] ;
wire \operand2[17] ;
wire \operand2[16] ;
wire \operand2[15] ;
wire \operand2[14] ;
wire \operand2[13] ;
wire \operand2[12] ;
wire \operand2[11] ;
wire \operand2[10] ;
wire \operand2[9] ;
wire \operand2[8] ;
wire \operand2[7] ;
wire \operand2[6] ;
wire \operand2[5] ;
wire \operand2[4] ;
wire \operand2[3] ;
wire \operand2[2] ;
wire \operand2[1] ;
wire \operand2[0] ;
wire \result[63] ;
wire \result[62] ;
wire \result[61] ;
wire \result[60] ;
wire \result[59] ;
wire \result[58] ;
wire \result[57] ;
wire \result[56] ;
wire \result[55] ;
wire \result[54] ;
wire \result[53] ;
wire \result[52] ;
wire \result[51] ;
wire \result[50] ;
wire \result[49] ;
wire \result[48] ;
wire \result[47] ;
wire \result[46] ;
wire \result[45] ;
wire \result[44] ;
wire \result[43] ;
wire \result[42] ;
wire \result[41] ;
wire \result[40] ;
wire \result[39] ;
wire \result[38] ;
wire \result[37] ;
wire \result[36] ;
wire \result[35] ;
wire \result[34] ;
wire \result[33] ;
wire \result[32] ;
wire \result[31] ;
wire \result[30] ;
wire \result[29] ;
wire \result[28] ;
wire \result[27] ;
wire \result[26] ;
wire \result[25] ;
wire \result[24] ;
wire \result[23] ;
wire \result[22] ;
wire \result[21] ;
wire \result[20] ;
wire \result[19] ;
wire \result[18] ;
wire \result[17] ;
wire \result[16] ;
wire \result[15] ;
wire \result[14] ;
wire \result[13] ;
wire \result[12] ;
wire \result[11] ;
wire \result[10] ;
wire \result[9] ;
wire \result[8] ;
wire \result[7] ;
wire \result[6] ;
wire \result[5] ;
wire \result[4] ;
wire \result[3] ;
wire \result[2] ;
wire \result[1] ;
wire \result[0] ;
wire CTS_n660;
wire CTS_n647;
wire CTS_n650;
wire CTS_n663;
wire CLOCK_n694;
wire CTS_n653;
wire CLOCK_slh__n955;
wire CLOCK_slh__n957;
wire CLOCK_slh__n959;
wire CLOCK_slh__n961;
wire CLOCK_slh__n963;
wire CLOCK_slh__n965;
wire CLOCK_slh__n967;
wire CLOCK_slh__n969;
wire CLOCK_slh__n971;
wire CLOCK_slh__n973;
wire CLOCK_slh__n975;
wire CLOCK_slh__n977;
wire CLOCK_slh__n979;
wire CLOCK_slh__n981;
wire CLOCK_slh__n983;
wire CLOCK_slh__n985;
wire CLOCK_slh__n987;
wire CLOCK_slh__n989;
wire CLOCK_slh__n991;
wire CLOCK_slh__n993;
wire CLOCK_slh__n995;
wire CLOCK_slh__n997;
wire CLOCK_slh__n999;
wire CLOCK_slh__n1001;
wire CLOCK_slh__n1003;
wire CLOCK_slh__n1005;
wire CLOCK_slh__n1007;
wire CLOCK_slh__n1009;
wire CLOCK_slh__n1011;
wire CLOCK_slh__n1013;
wire CLOCK_slh__n1015;
wire CLOCK_slh__n1017;
wire CLOCK_slh__n1019;
wire CLOCK_slh__n1021;
wire CLOCK_slh__n1023;
wire CLOCK_slh__n1025;
wire CLOCK_slh__n1027;
wire CLOCK_slh__n1029;
wire CLOCK_slh__n1031;
wire CLOCK_slh__n1033;
wire CLOCK_slh__n1035;
wire CLOCK_slh__n1037;
wire CLOCK_slh__n1039;
wire CLOCK_slh__n1041;
wire CLOCK_slh__n1043;
wire CLOCK_slh__n1045;
wire CLOCK_slh__n1047;
wire CLOCK_slh__n1049;
wire CLOCK_slh__n1051;
wire CLOCK_sph__n1055;
wire CLOCK_sph__n1057;


Register__parameterized0 Register_inst3 (.out ({out[63], out[62], out[61], out[60], 
    out[59], out[58], out[57], out[56], out[55], out[54], out[53], out[52], out[51], 
    out[50], out[49], out[48], out[47], out[46], out[45], out[44], out[43], out[42], 
    out[41], out[40], out[39], out[38], out[37], out[36], out[35], out[34], out[33], 
    out[32], out[31], out[30], out[29], out[28], out[27], out[26], out[25], out[24], 
    out[23], out[22], out[21], out[20], out[19], out[18], out[17], out[16], out[15], 
    out[14], out[13], out[12], out[11], out[10], out[9], out[8], out[7], out[6], 
    out[5], out[4], out[3], out[2], out[1], out[0]}), .clk_CTSPP_157 (CTS_n663), .in ({
    \result[63] , \result[62] , \result[61] , \result[60] , \result[59] , \result[58] , 
    \result[57] , \result[56] , \result[55] , \result[54] , \result[53] , \result[52] , 
    \result[51] , \result[50] , \result[49] , \result[48] , \result[47] , \result[46] , 
    \result[45] , \result[44] , \result[43] , \result[42] , \result[41] , \result[40] , 
    \result[39] , \result[38] , \result[37] , \result[36] , \result[35] , \result[34] , 
    \result[33] , \result[32] , \result[31] , \result[30] , \result[29] , \result[28] , 
    \result[27] , \result[26] , \result[25] , \result[24] , \result[23] , \result[22] , 
    \result[21] , \result[20] , \result[19] , \result[18] , \result[17] , \result[16] , 
    \result[15] , \result[14] , \result[13] , \result[12] , \result[11] , \result[10] , 
    \result[9] , \result[8] , \result[7] , \result[6] , \result[5] , \result[4] , 
    \result[3] , \result[2] , \result[1] , \result[0] }), .clk_CTSPP_154 (CTS_n650)
    , .clk_CTSPP_156 (CTS_n660), .clk_CTSPP_159 (CLOCK_n694));
sequential_multiplier sequential_multiplier_inst (.out ({\result[63] , \result[62] , 
    \result[61] , \result[60] , \result[59] , \result[58] , \result[57] , \result[56] , 
    \result[55] , \result[54] , \result[53] , \result[52] , \result[51] , \result[50] , 
    \result[49] , \result[48] , \result[47] , \result[46] , \result[45] , \result[44] , 
    \result[43] , \result[42] , \result[41] , \result[40] , \result[39] , \result[38] , 
    \result[37] , \result[36] , \result[35] , \result[34] , \result[33] , \result[32] , 
    \result[31] , \result[30] , \result[29] , \result[28] , \result[27] , \result[26] , 
    \result[25] , \result[24] , \result[23] , \result[22] , \result[21] , \result[20] , 
    \result[19] , \result[18] , \result[17] , \result[16] , \result[15] , \result[14] , 
    \result[13] , \result[12] , \result[11] , \result[10] , \result[9] , \result[8] , 
    \result[7] , \result[6] , \result[5] , \result[4] , \result[3] , \result[2] , 
    \result[1] , \result[0] }), .clk_CTSPP_233 (CTS_n660), .in1 ({\operand1[31] , 
    \operand1[30] , \operand1[29] , \operand1[28] , \operand1[27] , \operand1[26] , 
    \operand1[25] , \operand1[24] , \operand1[23] , \operand1[22] , \operand1[21] , 
    \operand1[20] , \operand1[19] , \operand1[18] , \operand1[17] , \operand1[16] , 
    \operand1[15] , \operand1[14] , \operand1[13] , \operand1[12] , \operand1[11] , 
    \operand1[10] , \operand1[9] , \operand1[8] , \operand1[7] , \operand1[6] , \operand1[5] , 
    \operand1[4] , \operand1[3] , \operand1[2] , \operand1[1] , \operand1[0] }), .in2 ({
    \operand2[31] , \operand2[30] , \operand2[29] , \operand2[28] , \operand2[27] , 
    \operand2[26] , \operand2[25] , \operand2[24] , \operand2[23] , \operand2[22] , 
    \operand2[21] , \operand2[20] , \operand2[19] , \operand2[18] , \operand2[17] , 
    \operand2[16] , \operand2[15] , \operand2[14] , \operand2[13] , \operand2[12] , 
    \operand2[11] , \operand2[10] , \operand2[9] , \operand2[8] , \operand2[7] , 
    \operand2[6] , \operand2[5] , \operand2[4] , \operand2[3] , \operand2[2] , \operand2[1] , 
    \operand2[0] }), .rst (rst), .clk_CTSPP_229 (CTS_n647), .clk_CTSPP_230 (CTS_n650)
    , .clk_CTSPP_231 (CTS_n653), .clk_CTSPP_234 (CTS_n663), .clk_CTSPP_236 (CLOCK_n694));
Register Register_inst2 (.out ({\operand2[31] , \operand2[30] , \operand2[29] , \operand2[28] , 
    \operand2[27] , \operand2[26] , \operand2[25] , \operand2[24] , \operand2[23] , 
    \operand2[22] , \operand2[21] , \operand2[20] , \operand2[19] , \operand2[18] , 
    \operand2[17] , \operand2[16] , \operand2[15] , \operand2[14] , \operand2[13] , 
    \operand2[12] , \operand2[11] , \operand2[10] , \operand2[9] , \operand2[8] , 
    \operand2[7] , \operand2[6] , \operand2[5] , \operand2[4] , \operand2[3] , \operand2[2] , 
    \operand2[1] , \operand2[0] }), .clk_CTSPP_119 (CTS_n647), .clk_CTSPP_120 (CTS_n653)
    , .in ({CLOCK_slh_n824, CLOCK_slh_n844, CLOCK_slh_n914, CLOCK_slh_n909, CLOCK_slh_n804, 
    CLOCK_slh_n754, CLOCK_slh_n799, CLOCK_slh_n889, CLOCK_slh_n794, CLOCK_slh_n789, 
    CLOCK_slh_n784, CLOCK_slh_n779, CLOCK_slh_n774, CLOCK_slh_n769, CLOCK_slh_n764, 
    CLOCK_slh_n759, CLOCK_slh_n744, CLOCK_slh_n749, CLOCK_slh_n739, CLOCK_slh_n734, 
    CLOCK_slh_n729, in2[10], in2[9], in2[8], in2[7], CLOCK_slh_n719, CLOCK_slh_n724, 
    CLOCK_slh_n709, CLOCK_slh_n714, CLOCK_slh_n809, CLOCK_slh_n884, CLOCK_slh_n864})
    , .clk_CTSPP_122 (CTS_n660), .clk_CTSPP_125 (CLOCK_n694));
Register__0_13 Register_inst1 (.out ({\operand1[31] , \operand1[30] , \operand1[29] , 
    \operand1[28] , \operand1[27] , \operand1[26] , \operand1[25] , \operand1[24] , 
    \operand1[23] , \operand1[22] , \operand1[21] , \operand1[20] , \operand1[19] , 
    \operand1[18] , \operand1[17] , \operand1[16] , \operand1[15] , \operand1[14] , 
    \operand1[13] , \operand1[12] , \operand1[11] , \operand1[10] , \operand1[9] , 
    \operand1[8] , \operand1[7] , \operand1[6] , \operand1[5] , \operand1[4] , \operand1[3] , 
    \operand1[2] , \operand1[1] , \operand1[0] }), .clk_CTSPP_192 (CTS_n650), .in ({
    CLOCK_slh_n869, CLOCK_slh_n944, CLOCK_slh_n939, CLOCK_slh_n949, CLOCK_slh_n934, 
    CLOCK_slh_n929, CLOCK_slh_n879, CLOCK_slh_n904, CLOCK_slh_n874, CLOCK_slh_n854, 
    CLOCK_slh_n899, CLOCK_slh_n894, CLOCK_slh_n849, CLOCK_slh_n839, CLOCK_slh_n859, 
    CLOCK_slh_n819, CLOCK_slh_n834, CLOCK_slh_n919, CLOCK_slh_n924, CLOCK_slh_n829, 
    CLOCK_slh_n814, in1[10], CLOCK_slh_n954, in1[8], in1[7], CLOCK_slh_n699, CLOCK_slh_n704, 
    in1[4], in1[3], in1[2], in1[1], in1[0]}), .clk_CTSPP_191 (CTS_n647), .clk_CTSPP_193 (CTS_n653)
    , .clk_CTSPP_195 (CTS_n660), .clk_CTSPP_196 (CTS_n663), .clk_CTSPP_198 (CLOCK_n694));
CLKBUF_X3 CTS_L1_c1_c27 (.Z (CLOCK_n694), .A (clk));
CLKBUF_X1 CLOCK_slh__c31 (.Z (CLOCK_slh__n1027), .A (in1[6]));
CLKBUF_X1 CLOCK_slh__c33 (.Z (CLOCK_slh__n1029), .A (in1[5]));
CLKBUF_X1 CLOCK_slh__c35 (.Z (CLOCK_slh__n981), .A (in2[4]));
CLKBUF_X1 CLOCK_slh__c37 (.Z (CLOCK_slh__n975), .A (in2[3]));
CLKBUF_X1 CLOCK_slh__c39 (.Z (CLOCK_slh__n977), .A (in2[6]));
CLKBUF_X1 CLOCK_slh__c41 (.Z (CLOCK_slh__n955), .A (in2[5]));
CLKBUF_X1 CLOCK_slh__c43 (.Z (CLOCK_slh__n1049), .A (in2[11]));
CLKBUF_X1 CLOCK_slh__c45 (.Z (CLOCK_slh__n957), .A (in2[12]));
CLKBUF_X1 CLOCK_slh__c47 (.Z (CLOCK_slh__n979), .A (in2[13]));
CLKBUF_X1 CLOCK_slh__c49 (.Z (CLOCK_slh__n959), .A (in2[15]));
CLKBUF_X1 CLOCK_slh__c51 (.Z (CLOCK_slh__n983), .A (in2[14]));
CLKBUF_X1 CLOCK_slh__c53 (.Z (CLOCK_slh__n961), .A (in2[26]));
CLKBUF_X1 CLOCK_slh__c55 (.Z (CLOCK_slh__n965), .A (in2[16]));
CLKBUF_X1 CLOCK_slh__c57 (.Z (CLOCK_slh__n1015), .A (in2[17]));
CLKBUF_X1 CLOCK_slh__c59 (.Z (CLOCK_slh__n967), .A (in2[18]));
CLKBUF_X1 CLOCK_slh__c61 (.Z (CLOCK_slh__n963), .A (in2[19]));
CLKBUF_X1 CLOCK_slh__c63 (.Z (CLOCK_slh__n969), .A (in2[20]));
CLKBUF_X1 CLOCK_slh__c65 (.Z (CLOCK_slh__n987), .A (in2[21]));
CLKBUF_X1 CLOCK_slh__c67 (.Z (CLOCK_slh__n973), .A (in2[22]));
CLKBUF_X1 CLOCK_slh__c69 (.Z (CLOCK_slh__n985), .A (in2[23]));
CLKBUF_X1 CLOCK_slh__c71 (.Z (CLOCK_slh__n1013), .A (in2[25]));
CLKBUF_X1 CLOCK_slh__c73 (.Z (CLOCK_slh__n1011), .A (in2[27]));
CLKBUF_X1 CLOCK_slh__c75 (.Z (CLOCK_slh__n971), .A (in2[2]));
CLKBUF_X1 CLOCK_slh__c77 (.Z (CLOCK_slh__n1003), .A (in1[11]));
CLKBUF_X1 CLOCK_slh__c79 (.Z (CLOCK_slh__n993), .A (in1[16]));
CLKBUF_X1 CLOCK_slh__c81 (.Z (CLOCK_slh__n989), .A (in2[31]));
CLKBUF_X1 CLOCK_slh__c83 (.Z (CLOCK_slh__n1005), .A (in1[12]));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_slh__n1019), .A (in1[15]));
CLKBUF_X1 CLOCK_slh__c87 (.Z (CLOCK_slh__n1017), .A (in1[18]));
CLKBUF_X1 CLOCK_slh__c89 (.Z (CLOCK_slh__n1031), .A (in2[30]));
CLKBUF_X1 CLOCK_slh__c91 (.Z (CLOCK_slh__n1023), .A (in1[19]));
CLKBUF_X1 CLOCK_slh__c93 (.Z (CLOCK_slh__n1021), .A (in1[22]));
CLKBUF_X1 CLOCK_slh__c95 (.Z (CLOCK_slh__n1007), .A (in1[17]));
CLKBUF_X1 CLOCK_slh__c97 (.Z (CLOCK_slh__n1009), .A (in2[0]));
CLKBUF_X1 CLOCK_slh__c99 (.Z (CLOCK_slh__n995), .A (in1[31]));
CLKBUF_X1 CLOCK_slh__c101 (.Z (CLOCK_slh__n1035), .A (in1[23]));
CLKBUF_X1 CLOCK_slh__c103 (.Z (CLOCK_slh__n1025), .A (in1[25]));
CLKBUF_X1 CLOCK_slh__c105 (.Z (CLOCK_slh__n991), .A (in2[1]));
CLKBUF_X1 CLOCK_slh__c107 (.Z (CLOCK_slh__n999), .A (in2[24]));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh__n1043), .A (in1[20]));
CLKBUF_X1 CLOCK_slh__c111 (.Z (CLOCK_slh__n997), .A (in1[21]));
CLKBUF_X1 CLOCK_slh__c113 (.Z (CLOCK_slh__n1045), .A (in1[24]));
CLKBUF_X1 CLOCK_slh__c115 (.Z (CLOCK_slh__n1033), .A (in2[28]));
CLKBUF_X1 CLOCK_slh__c117 (.Z (CLOCK_slh__n1001), .A (in2[29]));
CLKBUF_X1 CLOCK_slh__c119 (.Z (CLOCK_sph__n1055), .A (in1[14]));
CLKBUF_X1 CLOCK_slh__c121 (.Z (CLOCK_slh__n1039), .A (in1[13]));
CLKBUF_X1 CLOCK_slh__c123 (.Z (CLOCK_slh__n1037), .A (in1[26]));
CLKBUF_X1 CLOCK_slh__c125 (.Z (CLOCK_slh__n1041), .A (in1[27]));
CLKBUF_X1 CLOCK_slh__c127 (.Z (CLOCK_slh__n1047), .A (in1[29]));
CLKBUF_X1 CLOCK_slh__c129 (.Z (CLOCK_sph__n1057), .A (in1[30]));
CLKBUF_X1 CLOCK_slh__c131 (.Z (CLOCK_slh__n1051), .A (in1[28]));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_slh_n954), .A (in1[9]));
CLKBUF_X1 CLOCK_slh__c135 (.Z (CLOCK_slh_n724), .A (CLOCK_slh__n955));
CLKBUF_X1 CLOCK_slh__c137 (.Z (CLOCK_slh_n734), .A (CLOCK_slh__n957));
CLKBUF_X1 CLOCK_slh__c139 (.Z (CLOCK_slh_n744), .A (CLOCK_slh__n959));
CLKBUF_X1 CLOCK_slh__c141 (.Z (CLOCK_slh_n754), .A (CLOCK_slh__n961));
CLKBUF_X1 CLOCK_slh__c143 (.Z (CLOCK_slh_n774), .A (CLOCK_slh__n963));
CLKBUF_X1 CLOCK_slh__c145 (.Z (CLOCK_slh_n759), .A (CLOCK_slh__n965));
CLKBUF_X1 CLOCK_slh__c147 (.Z (CLOCK_slh_n769), .A (CLOCK_slh__n967));
CLKBUF_X1 CLOCK_slh__c149 (.Z (CLOCK_slh_n779), .A (CLOCK_slh__n969));
CLKBUF_X1 CLOCK_slh__c151 (.Z (CLOCK_slh_n809), .A (CLOCK_slh__n971));
CLKBUF_X1 CLOCK_slh__c153 (.Z (CLOCK_slh_n789), .A (CLOCK_slh__n973));
CLKBUF_X1 CLOCK_slh__c155 (.Z (CLOCK_slh_n714), .A (CLOCK_slh__n975));
CLKBUF_X1 CLOCK_slh__c157 (.Z (CLOCK_slh_n719), .A (CLOCK_slh__n977));
CLKBUF_X1 CLOCK_slh__c159 (.Z (CLOCK_slh_n739), .A (CLOCK_slh__n979));
CLKBUF_X1 CLOCK_slh__c161 (.Z (CLOCK_slh_n709), .A (CLOCK_slh__n981));
CLKBUF_X1 CLOCK_slh__c163 (.Z (CLOCK_slh_n749), .A (CLOCK_slh__n983));
CLKBUF_X1 CLOCK_slh__c165 (.Z (CLOCK_slh_n794), .A (CLOCK_slh__n985));
CLKBUF_X1 CLOCK_slh__c167 (.Z (CLOCK_slh_n784), .A (CLOCK_slh__n987));
CLKBUF_X1 CLOCK_slh__c169 (.Z (CLOCK_slh_n824), .A (CLOCK_slh__n989));
CLKBUF_X1 CLOCK_slh__c171 (.Z (CLOCK_slh_n884), .A (CLOCK_slh__n991));
CLKBUF_X1 CLOCK_slh__c173 (.Z (CLOCK_slh_n819), .A (CLOCK_slh__n993));
CLKBUF_X1 CLOCK_slh__c175 (.Z (CLOCK_slh_n869), .A (CLOCK_slh__n995));
CLKBUF_X1 CLOCK_slh__c177 (.Z (CLOCK_slh_n899), .A (CLOCK_slh__n997));
CLKBUF_X1 CLOCK_slh__c179 (.Z (CLOCK_slh_n889), .A (CLOCK_slh__n999));
CLKBUF_X1 CLOCK_slh__c181 (.Z (CLOCK_slh_n914), .A (CLOCK_slh__n1001));
CLKBUF_X1 CLOCK_slh__c183 (.Z (CLOCK_slh_n814), .A (CLOCK_slh__n1003));
CLKBUF_X1 CLOCK_slh__c185 (.Z (CLOCK_slh_n829), .A (CLOCK_slh__n1005));
CLKBUF_X1 CLOCK_slh__c187 (.Z (CLOCK_slh_n859), .A (CLOCK_slh__n1007));
CLKBUF_X1 CLOCK_slh__c189 (.Z (CLOCK_slh_n864), .A (CLOCK_slh__n1009));
CLKBUF_X1 CLOCK_slh__c191 (.Z (CLOCK_slh_n804), .A (CLOCK_slh__n1011));
CLKBUF_X1 CLOCK_slh__c193 (.Z (CLOCK_slh_n799), .A (CLOCK_slh__n1013));
CLKBUF_X1 CLOCK_slh__c195 (.Z (CLOCK_slh_n764), .A (CLOCK_slh__n1015));
CLKBUF_X1 CLOCK_slh__c197 (.Z (CLOCK_slh_n839), .A (CLOCK_slh__n1017));
CLKBUF_X1 CLOCK_slh__c199 (.Z (CLOCK_slh_n834), .A (CLOCK_slh__n1019));
CLKBUF_X1 CLOCK_slh__c201 (.Z (CLOCK_slh_n854), .A (CLOCK_slh__n1021));
CLKBUF_X1 CLOCK_slh__c203 (.Z (CLOCK_slh_n849), .A (CLOCK_slh__n1023));
CLKBUF_X1 CLOCK_slh__c205 (.Z (CLOCK_slh_n879), .A (CLOCK_slh__n1025));
CLKBUF_X1 CLOCK_slh__c207 (.Z (CLOCK_slh_n699), .A (CLOCK_slh__n1027));
CLKBUF_X1 CLOCK_slh__c209 (.Z (CLOCK_slh_n704), .A (CLOCK_slh__n1029));
CLKBUF_X1 CLOCK_slh__c211 (.Z (CLOCK_slh_n844), .A (CLOCK_slh__n1031));
CLKBUF_X1 CLOCK_slh__c213 (.Z (CLOCK_slh_n909), .A (CLOCK_slh__n1033));
CLKBUF_X1 CLOCK_slh__c215 (.Z (CLOCK_slh_n874), .A (CLOCK_slh__n1035));
CLKBUF_X1 CLOCK_slh__c217 (.Z (CLOCK_slh_n929), .A (CLOCK_slh__n1037));
CLKBUF_X1 CLOCK_slh__c219 (.Z (CLOCK_slh_n924), .A (CLOCK_slh__n1039));
CLKBUF_X1 CLOCK_slh__c221 (.Z (CLOCK_slh_n934), .A (CLOCK_slh__n1041));
CLKBUF_X1 CLOCK_slh__c223 (.Z (CLOCK_slh_n894), .A (CLOCK_slh__n1043));
CLKBUF_X1 CLOCK_slh__c225 (.Z (CLOCK_slh_n904), .A (CLOCK_slh__n1045));
CLKBUF_X1 CLOCK_slh__c227 (.Z (CLOCK_slh_n939), .A (CLOCK_slh__n1047));
CLKBUF_X1 CLOCK_slh__c229 (.Z (CLOCK_slh_n729), .A (CLOCK_slh__n1049));
CLKBUF_X1 CLOCK_slh__c231 (.Z (CLOCK_slh_n949), .A (CLOCK_slh__n1051));
CLKBUF_X1 CLOCK_sph__c235 (.Z (CLOCK_slh_n919), .A (CLOCK_sph__n1055));
CLKBUF_X1 CLOCK_sph__c237 (.Z (CLOCK_slh_n944), .A (CLOCK_sph__n1057));

endmodule //SequentialMultiplierIntegerated


