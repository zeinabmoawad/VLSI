/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Dec 15 00:06:12 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1754676415 */

module datapath__0_130(p_0, p_1, p_2, p_3, p_4, p_5, p_6, p_7, p_8, p_9, p_10, 
      p_11, p_12, p_13, p_14, p_15, p_16, p_17, p_18, p_19, p_20, p_21, p_22, 
      p_23, p_24, p_25, p_26, p_27, p_28, p_29, p_30, out, out31);
   input [63:0]p_0;
   input [63:0]p_1;
   input [63:0]p_2;
   input [63:0]p_3;
   input [63:0]p_4;
   input [63:0]p_5;
   input [63:0]p_6;
   input [63:0]p_7;
   input [63:0]p_8;
   input [63:0]p_9;
   input [63:0]p_10;
   input [63:0]p_11;
   input [63:0]p_12;
   input [63:0]p_13;
   input [63:0]p_14;
   input [63:0]p_15;
   input [63:0]p_16;
   input [63:0]p_17;
   input [63:0]p_18;
   input [63:0]p_19;
   input [63:0]p_20;
   input [63:0]p_21;
   input [63:0]p_22;
   input [63:0]p_23;
   input [63:0]p_24;
   input [63:0]p_25;
   input [63:0]p_26;
   input [63:0]p_27;
   input [63:0]p_28;
   input [63:0]p_29;
   input [63:0]p_30;
   input [63:0]out;
   output [63:0]out31;

   HA_X1 i_0 (.A(p_0[2]), .B(p_1[2]), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(p_0[3]), .B(p_1[3]), .CI(p_2[3]), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(out[3]), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(p_2[4]), .CO(n_7), .S(n_6));
   FA_X1 i_4 (.A(p_3[4]), .B(out[4]), .CI(n_5), .CO(n_9), .S(n_8));
   HA_X1 i_5 (.A(n_3), .B(n_8), .CO(n_11), .S(n_10));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(p_2[5]), .CO(n_13), .S(n_12));
   FA_X1 i_7 (.A(p_3[5]), .B(p_4[5]), .CI(out[5]), .CO(n_15), .S(n_14));
   FA_X1 i_8 (.A(n_7), .B(n_9), .CI(n_14), .CO(n_17), .S(n_16));
   HA_X1 i_9 (.A(n_12), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_10 (.A(p_0[6]), .B(p_1[6]), .CI(p_2[6]), .CO(n_21), .S(n_20));
   FA_X1 i_11 (.A(p_3[6]), .B(p_4[6]), .CI(p_5[6]), .CO(n_23), .S(n_22));
   FA_X1 i_12 (.A(out[6]), .B(n_15), .CI(n_13), .CO(n_25), .S(n_24));
   FA_X1 i_13 (.A(n_22), .B(n_20), .CI(n_24), .CO(n_27), .S(n_26));
   HA_X1 i_14 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_15 (.A(p_0[7]), .B(p_1[7]), .CI(p_2[7]), .CO(n_31), .S(n_30));
   FA_X1 i_16 (.A(p_3[7]), .B(p_4[7]), .CI(p_5[7]), .CO(n_33), .S(n_32));
   FA_X1 i_17 (.A(p_6[7]), .B(out[7]), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_18 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_19 (.A(n_32), .B(n_30), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_20 (.A(n_36), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_21 (.A(p_0[8]), .B(p_1[8]), .CI(p_2[8]), .CO(n_43), .S(n_42));
   FA_X1 i_22 (.A(p_3[8]), .B(p_4[8]), .CI(p_5[8]), .CO(n_45), .S(n_44));
   FA_X1 i_23 (.A(p_6[8]), .B(p_7[8]), .CI(out[8]), .CO(n_47), .S(n_46));
   FA_X1 i_24 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_48));
   FA_X1 i_25 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_51), .S(n_50));
   FA_X1 i_26 (.A(n_48), .B(n_37), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_27 (.A(n_39), .B(n_50), .CO(n_55), .S(n_54));
   FA_X1 i_28 (.A(p_0[9]), .B(p_1[9]), .CI(p_2[9]), .CO(n_57), .S(n_56));
   FA_X1 i_29 (.A(p_3[9]), .B(p_4[9]), .CI(p_5[9]), .CO(n_59), .S(n_58));
   FA_X1 i_30 (.A(p_6[9]), .B(p_7[9]), .CI(p_8[9]), .CO(n_61), .S(n_60));
   FA_X1 i_31 (.A(out[9]), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_32 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_64));
   FA_X1 i_33 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_67), .S(n_66));
   FA_X1 i_34 (.A(n_51), .B(n_64), .CI(n_66), .CO(n_69), .S(n_68));
   HA_X1 i_35 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_36 (.A(p_0[10]), .B(p_1[10]), .CI(p_2[10]), .CO(n_73), .S(n_72));
   FA_X1 i_37 (.A(p_3[10]), .B(p_4[10]), .CI(p_5[10]), .CO(n_75), .S(n_74));
   FA_X1 i_38 (.A(p_6[10]), .B(p_7[10]), .CI(p_8[10]), .CO(n_77), .S(n_76));
   FA_X1 i_39 (.A(p_9[10]), .B(out[10]), .CI(n_61), .CO(n_79), .S(n_78));
   FA_X1 i_40 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_81), .S(n_80));
   FA_X1 i_41 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_83), .S(n_82));
   FA_X1 i_42 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_85), .S(n_84));
   FA_X1 i_43 (.A(n_67), .B(n_82), .CI(n_84), .CO(n_87), .S(n_86));
   HA_X1 i_44 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_45 (.A(p_0[11]), .B(p_1[11]), .CI(p_2[11]), .CO(n_91), .S(n_90));
   FA_X1 i_46 (.A(p_3[11]), .B(p_4[11]), .CI(p_5[11]), .CO(n_93), .S(n_92));
   FA_X1 i_47 (.A(p_6[11]), .B(p_7[11]), .CI(p_8[11]), .CO(n_95), .S(n_94));
   FA_X1 i_48 (.A(p_9[11]), .B(p_10[11]), .CI(out[11]), .CO(n_97), .S(n_96));
   FA_X1 i_49 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_99), .S(n_98));
   FA_X1 i_50 (.A(n_79), .B(n_96), .CI(n_94), .CO(n_101), .S(n_100));
   FA_X1 i_51 (.A(n_92), .B(n_90), .CI(n_81), .CO(n_103), .S(n_102));
   FA_X1 i_52 (.A(n_98), .B(n_83), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_53 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_54 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   FA_X1 i_55 (.A(p_0[12]), .B(p_1[12]), .CI(p_2[12]), .CO(n_111), .S(n_110));
   FA_X1 i_56 (.A(p_3[12]), .B(p_4[12]), .CI(p_5[12]), .CO(n_113), .S(n_112));
   FA_X1 i_57 (.A(p_6[12]), .B(p_7[12]), .CI(p_8[12]), .CO(n_115), .S(n_114));
   FA_X1 i_58 (.A(p_9[12]), .B(p_10[12]), .CI(p_11[12]), .CO(n_117), .S(n_116));
   FA_X1 i_59 (.A(out[12]), .B(n_97), .CI(n_95), .CO(n_119), .S(n_118));
   FA_X1 i_60 (.A(n_93), .B(n_91), .CI(n_99), .CO(n_121), .S(n_120));
   FA_X1 i_61 (.A(n_116), .B(n_114), .CI(n_112), .CO(n_123), .S(n_122));
   FA_X1 i_62 (.A(n_110), .B(n_120), .CI(n_118), .CO(n_125), .S(n_124));
   FA_X1 i_63 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_64 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   HA_X1 i_65 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_66 (.A(p_0[13]), .B(p_1[13]), .CI(p_2[13]), .CO(n_133), .S(n_132));
   FA_X1 i_67 (.A(p_3[13]), .B(p_4[13]), .CI(p_5[13]), .CO(n_135), .S(n_134));
   FA_X1 i_68 (.A(p_6[13]), .B(p_7[13]), .CI(p_8[13]), .CO(n_137), .S(n_136));
   FA_X1 i_69 (.A(p_9[13]), .B(p_10[13]), .CI(p_11[13]), .CO(n_139), .S(n_138));
   FA_X1 i_70 (.A(p_12[13]), .B(out[13]), .CI(n_117), .CO(n_141), .S(n_140));
   FA_X1 i_71 (.A(n_115), .B(n_113), .CI(n_111), .CO(n_143), .S(n_142));
   FA_X1 i_72 (.A(n_119), .B(n_140), .CI(n_138), .CO(n_145), .S(n_144));
   FA_X1 i_73 (.A(n_136), .B(n_134), .CI(n_132), .CO(n_147), .S(n_146));
   FA_X1 i_74 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_75 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_76 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_77 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   FA_X1 i_78 (.A(p_0[14]), .B(p_1[14]), .CI(p_2[14]), .CO(n_157), .S(n_156));
   FA_X1 i_79 (.A(p_3[14]), .B(p_4[14]), .CI(p_5[14]), .CO(n_159), .S(n_158));
   FA_X1 i_80 (.A(p_6[14]), .B(p_7[14]), .CI(p_8[14]), .CO(n_161), .S(n_160));
   FA_X1 i_81 (.A(p_9[14]), .B(p_10[14]), .CI(p_11[14]), .CO(n_163), .S(n_162));
   FA_X1 i_82 (.A(p_12[14]), .B(p_13[14]), .CI(out[14]), .CO(n_165), .S(n_164));
   FA_X1 i_83 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_167), .S(n_166));
   FA_X1 i_84 (.A(n_133), .B(n_143), .CI(n_141), .CO(n_169), .S(n_168));
   FA_X1 i_85 (.A(n_164), .B(n_162), .CI(n_160), .CO(n_171), .S(n_170));
   FA_X1 i_86 (.A(n_158), .B(n_156), .CI(n_166), .CO(n_173), .S(n_172));
   FA_X1 i_87 (.A(n_147), .B(n_145), .CI(n_168), .CO(n_175), .S(n_174));
   FA_X1 i_88 (.A(n_149), .B(n_172), .CI(n_170), .CO(n_177), .S(n_176));
   FA_X1 i_89 (.A(n_174), .B(n_151), .CI(n_176), .CO(n_179), .S(n_178));
   HA_X1 i_90 (.A(n_153), .B(n_155), .CO(n_181), .S(n_180));
   FA_X1 i_91 (.A(p_0[15]), .B(p_1[15]), .CI(p_2[15]), .CO(n_183), .S(n_182));
   FA_X1 i_92 (.A(p_3[15]), .B(p_4[15]), .CI(p_5[15]), .CO(n_185), .S(n_184));
   FA_X1 i_93 (.A(p_6[15]), .B(p_7[15]), .CI(p_8[15]), .CO(n_187), .S(n_186));
   FA_X1 i_94 (.A(p_9[15]), .B(p_10[15]), .CI(p_11[15]), .CO(n_189), .S(n_188));
   FA_X1 i_95 (.A(p_12[15]), .B(p_13[15]), .CI(p_14[15]), .CO(n_191), .S(n_190));
   FA_X1 i_96 (.A(out[15]), .B(n_165), .CI(n_163), .CO(n_193), .S(n_192));
   FA_X1 i_97 (.A(n_161), .B(n_159), .CI(n_157), .CO(n_195), .S(n_194));
   FA_X1 i_98 (.A(n_167), .B(n_190), .CI(n_188), .CO(n_197), .S(n_196));
   FA_X1 i_99 (.A(n_186), .B(n_184), .CI(n_182), .CO(n_199), .S(n_198));
   FA_X1 i_100 (.A(n_169), .B(n_194), .CI(n_192), .CO(n_201), .S(n_200));
   FA_X1 i_101 (.A(n_171), .B(n_173), .CI(n_198), .CO(n_203), .S(n_202));
   FA_X1 i_102 (.A(n_196), .B(n_175), .CI(n_200), .CO(n_205), .S(n_204));
   FA_X1 i_103 (.A(n_177), .B(n_202), .CI(n_204), .CO(n_207), .S(n_206));
   HA_X1 i_104 (.A(n_179), .B(n_181), .CO(n_209), .S(n_208));
   FA_X1 i_105 (.A(p_0[16]), .B(p_1[16]), .CI(p_2[16]), .CO(n_211), .S(n_210));
   FA_X1 i_106 (.A(p_3[16]), .B(p_4[16]), .CI(p_5[16]), .CO(n_213), .S(n_212));
   FA_X1 i_107 (.A(p_6[16]), .B(p_7[16]), .CI(p_8[16]), .CO(n_215), .S(n_214));
   FA_X1 i_108 (.A(p_9[16]), .B(p_10[16]), .CI(p_11[16]), .CO(n_217), .S(n_216));
   FA_X1 i_109 (.A(p_12[16]), .B(p_13[16]), .CI(p_14[16]), .CO(n_219), .S(n_218));
   FA_X1 i_110 (.A(p_15[16]), .B(out[16]), .CI(n_191), .CO(n_221), .S(n_220));
   FA_X1 i_111 (.A(n_189), .B(n_187), .CI(n_185), .CO(n_223), .S(n_222));
   FA_X1 i_112 (.A(n_183), .B(n_195), .CI(n_193), .CO(n_225), .S(n_224));
   FA_X1 i_113 (.A(n_220), .B(n_218), .CI(n_216), .CO(n_227), .S(n_226));
   FA_X1 i_114 (.A(n_214), .B(n_212), .CI(n_210), .CO(n_229), .S(n_228));
   FA_X1 i_115 (.A(n_222), .B(n_199), .CI(n_197), .CO(n_231), .S(n_230));
   FA_X1 i_116 (.A(n_224), .B(n_201), .CI(n_228), .CO(n_233), .S(n_232));
   FA_X1 i_117 (.A(n_226), .B(n_230), .CI(n_203), .CO(n_235), .S(n_234));
   FA_X1 i_118 (.A(n_232), .B(n_205), .CI(n_234), .CO(n_237), .S(n_236));
   HA_X1 i_119 (.A(n_207), .B(n_209), .CO(n_239), .S(n_238));
   FA_X1 i_120 (.A(p_0[17]), .B(p_1[17]), .CI(p_2[17]), .CO(n_241), .S(n_240));
   FA_X1 i_121 (.A(p_3[17]), .B(p_4[17]), .CI(p_5[17]), .CO(n_243), .S(n_242));
   FA_X1 i_122 (.A(p_6[17]), .B(p_7[17]), .CI(p_8[17]), .CO(n_245), .S(n_244));
   FA_X1 i_123 (.A(p_9[17]), .B(p_10[17]), .CI(p_11[17]), .CO(n_247), .S(n_246));
   FA_X1 i_124 (.A(p_12[17]), .B(p_13[17]), .CI(p_14[17]), .CO(n_249), .S(n_248));
   FA_X1 i_125 (.A(p_15[17]), .B(p_16[17]), .CI(out[17]), .CO(n_251), .S(n_250));
   FA_X1 i_126 (.A(n_219), .B(n_217), .CI(n_215), .CO(n_253), .S(n_252));
   FA_X1 i_127 (.A(n_213), .B(n_211), .CI(n_223), .CO(n_255), .S(n_254));
   FA_X1 i_128 (.A(n_221), .B(n_250), .CI(n_248), .CO(n_257), .S(n_256));
   FA_X1 i_129 (.A(n_246), .B(n_244), .CI(n_242), .CO(n_259), .S(n_258));
   FA_X1 i_130 (.A(n_240), .B(n_225), .CI(n_254), .CO(n_261), .S(n_260));
   FA_X1 i_131 (.A(n_252), .B(n_229), .CI(n_227), .CO(n_263), .S(n_262));
   FA_X1 i_132 (.A(n_231), .B(n_258), .CI(n_256), .CO(n_265), .S(n_264));
   FA_X1 i_133 (.A(n_260), .B(n_262), .CI(n_233), .CO(n_267), .S(n_266));
   FA_X1 i_134 (.A(n_235), .B(n_264), .CI(n_266), .CO(n_269), .S(n_268));
   HA_X1 i_135 (.A(n_237), .B(n_239), .CO(n_271), .S(n_270));
   FA_X1 i_136 (.A(p_0[18]), .B(p_1[18]), .CI(p_2[18]), .CO(n_273), .S(n_272));
   FA_X1 i_137 (.A(p_3[18]), .B(p_4[18]), .CI(p_5[18]), .CO(n_275), .S(n_274));
   FA_X1 i_138 (.A(p_6[18]), .B(p_7[18]), .CI(p_8[18]), .CO(n_277), .S(n_276));
   FA_X1 i_139 (.A(p_9[18]), .B(p_10[18]), .CI(p_11[18]), .CO(n_279), .S(n_278));
   FA_X1 i_140 (.A(p_12[18]), .B(p_13[18]), .CI(p_14[18]), .CO(n_281), .S(n_280));
   FA_X1 i_141 (.A(p_15[18]), .B(p_16[18]), .CI(p_17[18]), .CO(n_283), .S(n_282));
   FA_X1 i_142 (.A(out[18]), .B(n_251), .CI(n_249), .CO(n_285), .S(n_284));
   FA_X1 i_143 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_287), .S(n_286));
   FA_X1 i_144 (.A(n_241), .B(n_253), .CI(n_282), .CO(n_289), .S(n_288));
   FA_X1 i_145 (.A(n_280), .B(n_278), .CI(n_276), .CO(n_291), .S(n_290));
   FA_X1 i_146 (.A(n_274), .B(n_272), .CI(n_255), .CO(n_293), .S(n_292));
   FA_X1 i_147 (.A(n_286), .B(n_284), .CI(n_259), .CO(n_295), .S(n_294));
   FA_X1 i_148 (.A(n_257), .B(n_288), .CI(n_263), .CO(n_297), .S(n_296));
   FA_X1 i_149 (.A(n_261), .B(n_292), .CI(n_290), .CO(n_299), .S(n_298));
   FA_X1 i_150 (.A(n_294), .B(n_265), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_151 (.A(n_267), .B(n_298), .CI(n_300), .CO(n_303), .S(n_302));
   HA_X1 i_152 (.A(n_269), .B(n_302), .CO(n_305), .S(n_304));
   FA_X1 i_153 (.A(p_0[19]), .B(p_1[19]), .CI(p_2[19]), .CO(n_307), .S(n_306));
   FA_X1 i_154 (.A(p_3[19]), .B(p_4[19]), .CI(p_5[19]), .CO(n_309), .S(n_308));
   FA_X1 i_155 (.A(p_6[19]), .B(p_7[19]), .CI(p_8[19]), .CO(n_311), .S(n_310));
   FA_X1 i_156 (.A(p_9[19]), .B(p_10[19]), .CI(p_11[19]), .CO(n_313), .S(n_312));
   FA_X1 i_157 (.A(p_12[19]), .B(p_13[19]), .CI(p_14[19]), .CO(n_315), .S(n_314));
   FA_X1 i_158 (.A(p_15[19]), .B(p_16[19]), .CI(p_17[19]), .CO(n_317), .S(n_316));
   FA_X1 i_159 (.A(p_18[19]), .B(out[19]), .CI(n_283), .CO(n_319), .S(n_318));
   FA_X1 i_160 (.A(n_281), .B(n_279), .CI(n_277), .CO(n_321), .S(n_320));
   FA_X1 i_161 (.A(n_275), .B(n_273), .CI(n_287), .CO(n_323), .S(n_322));
   FA_X1 i_162 (.A(n_285), .B(n_318), .CI(n_316), .CO(n_325), .S(n_324));
   FA_X1 i_163 (.A(n_314), .B(n_312), .CI(n_310), .CO(n_327), .S(n_326));
   FA_X1 i_164 (.A(n_308), .B(n_306), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_165 (.A(n_320), .B(n_291), .CI(n_289), .CO(n_331), .S(n_330));
   FA_X1 i_166 (.A(n_293), .B(n_295), .CI(n_328), .CO(n_333), .S(n_332));
   FA_X1 i_167 (.A(n_326), .B(n_324), .CI(n_297), .CO(n_335), .S(n_334));
   FA_X1 i_168 (.A(n_330), .B(n_299), .CI(n_332), .CO(n_337), .S(n_336));
   FA_X1 i_169 (.A(n_334), .B(n_301), .CI(n_336), .CO(n_339), .S(n_338));
   HA_X1 i_170 (.A(n_303), .B(n_338), .CO(n_341), .S(n_340));
   FA_X1 i_171 (.A(p_0[20]), .B(p_1[20]), .CI(p_2[20]), .CO(n_343), .S(n_342));
   FA_X1 i_172 (.A(p_3[20]), .B(p_4[20]), .CI(p_5[20]), .CO(n_345), .S(n_344));
   FA_X1 i_173 (.A(p_6[20]), .B(p_7[20]), .CI(p_8[20]), .CO(n_347), .S(n_346));
   FA_X1 i_174 (.A(p_9[20]), .B(p_10[20]), .CI(p_11[20]), .CO(n_349), .S(n_348));
   FA_X1 i_175 (.A(p_12[20]), .B(p_13[20]), .CI(p_14[20]), .CO(n_351), .S(n_350));
   FA_X1 i_176 (.A(p_15[20]), .B(p_16[20]), .CI(p_17[20]), .CO(n_353), .S(n_352));
   FA_X1 i_177 (.A(p_18[20]), .B(p_19[20]), .CI(out[20]), .CO(n_355), .S(n_354));
   FA_X1 i_178 (.A(n_317), .B(n_315), .CI(n_313), .CO(n_357), .S(n_356));
   FA_X1 i_179 (.A(n_311), .B(n_309), .CI(n_307), .CO(n_359), .S(n_358));
   FA_X1 i_180 (.A(n_321), .B(n_319), .CI(n_354), .CO(n_361), .S(n_360));
   FA_X1 i_181 (.A(n_352), .B(n_350), .CI(n_348), .CO(n_363), .S(n_362));
   FA_X1 i_182 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_365), .S(n_364));
   FA_X1 i_183 (.A(n_323), .B(n_358), .CI(n_356), .CO(n_367), .S(n_366));
   FA_X1 i_184 (.A(n_327), .B(n_325), .CI(n_360), .CO(n_369), .S(n_368));
   FA_X1 i_185 (.A(n_331), .B(n_329), .CI(n_364), .CO(n_371), .S(n_370));
   FA_X1 i_186 (.A(n_362), .B(n_368), .CI(n_366), .CO(n_373), .S(n_372));
   FA_X1 i_187 (.A(n_333), .B(n_335), .CI(n_370), .CO(n_375), .S(n_374));
   FA_X1 i_188 (.A(n_337), .B(n_372), .CI(n_374), .CO(n_377), .S(n_376));
   HA_X1 i_189 (.A(n_339), .B(n_341), .CO(n_379), .S(n_378));
   FA_X1 i_190 (.A(p_0[21]), .B(p_1[21]), .CI(p_2[21]), .CO(n_381), .S(n_380));
   FA_X1 i_191 (.A(p_3[21]), .B(p_4[21]), .CI(p_5[21]), .CO(n_383), .S(n_382));
   FA_X1 i_192 (.A(p_6[21]), .B(p_7[21]), .CI(p_8[21]), .CO(n_385), .S(n_384));
   FA_X1 i_193 (.A(p_9[21]), .B(p_10[21]), .CI(p_11[21]), .CO(n_387), .S(n_386));
   FA_X1 i_194 (.A(p_12[21]), .B(p_13[21]), .CI(p_14[21]), .CO(n_389), .S(n_388));
   FA_X1 i_195 (.A(p_15[21]), .B(p_16[21]), .CI(p_17[21]), .CO(n_391), .S(n_390));
   FA_X1 i_196 (.A(p_18[21]), .B(p_19[21]), .CI(p_20[21]), .CO(n_393), .S(n_392));
   FA_X1 i_197 (.A(out[21]), .B(n_355), .CI(n_353), .CO(n_395), .S(n_394));
   FA_X1 i_198 (.A(n_351), .B(n_349), .CI(n_347), .CO(n_397), .S(n_396));
   FA_X1 i_199 (.A(n_345), .B(n_343), .CI(n_359), .CO(n_399), .S(n_398));
   FA_X1 i_200 (.A(n_357), .B(n_392), .CI(n_390), .CO(n_401), .S(n_400));
   FA_X1 i_201 (.A(n_388), .B(n_386), .CI(n_384), .CO(n_403), .S(n_402));
   FA_X1 i_202 (.A(n_382), .B(n_380), .CI(n_398), .CO(n_405), .S(n_404));
   FA_X1 i_203 (.A(n_396), .B(n_394), .CI(n_365), .CO(n_407), .S(n_406));
   FA_X1 i_204 (.A(n_363), .B(n_361), .CI(n_367), .CO(n_409), .S(n_408));
   FA_X1 i_205 (.A(n_404), .B(n_402), .CI(n_400), .CO(n_411), .S(n_410));
   FA_X1 i_206 (.A(n_369), .B(n_408), .CI(n_406), .CO(n_413), .S(n_412));
   FA_X1 i_207 (.A(n_371), .B(n_373), .CI(n_410), .CO(n_415), .S(n_414));
   FA_X1 i_208 (.A(n_375), .B(n_412), .CI(n_414), .CO(n_417), .S(n_416));
   HA_X1 i_209 (.A(n_377), .B(n_416), .CO(n_419), .S(n_418));
   FA_X1 i_210 (.A(p_0[22]), .B(p_1[22]), .CI(p_2[22]), .CO(n_421), .S(n_420));
   FA_X1 i_211 (.A(p_3[22]), .B(p_4[22]), .CI(p_5[22]), .CO(n_423), .S(n_422));
   FA_X1 i_212 (.A(p_6[22]), .B(p_7[22]), .CI(p_8[22]), .CO(n_425), .S(n_424));
   FA_X1 i_213 (.A(p_9[22]), .B(p_10[22]), .CI(p_11[22]), .CO(n_427), .S(n_426));
   FA_X1 i_214 (.A(p_12[22]), .B(p_13[22]), .CI(p_14[22]), .CO(n_429), .S(n_428));
   FA_X1 i_215 (.A(p_15[22]), .B(p_16[22]), .CI(p_17[22]), .CO(n_431), .S(n_430));
   FA_X1 i_216 (.A(p_18[22]), .B(p_19[22]), .CI(p_20[22]), .CO(n_433), .S(n_432));
   FA_X1 i_217 (.A(p_21[22]), .B(out[22]), .CI(n_393), .CO(n_435), .S(n_434));
   FA_X1 i_218 (.A(n_391), .B(n_389), .CI(n_387), .CO(n_437), .S(n_436));
   FA_X1 i_219 (.A(n_385), .B(n_383), .CI(n_381), .CO(n_439), .S(n_438));
   FA_X1 i_220 (.A(n_397), .B(n_395), .CI(n_434), .CO(n_441), .S(n_440));
   FA_X1 i_221 (.A(n_432), .B(n_430), .CI(n_428), .CO(n_443), .S(n_442));
   FA_X1 i_222 (.A(n_426), .B(n_424), .CI(n_422), .CO(n_445), .S(n_444));
   FA_X1 i_223 (.A(n_420), .B(n_399), .CI(n_438), .CO(n_447), .S(n_446));
   FA_X1 i_224 (.A(n_436), .B(n_403), .CI(n_401), .CO(n_449), .S(n_448));
   FA_X1 i_225 (.A(n_440), .B(n_407), .CI(n_405), .CO(n_451), .S(n_450));
   FA_X1 i_226 (.A(n_444), .B(n_442), .CI(n_446), .CO(n_453), .S(n_452));
   FA_X1 i_227 (.A(n_409), .B(n_448), .CI(n_411), .CO(n_455), .S(n_454));
   FA_X1 i_228 (.A(n_450), .B(n_413), .CI(n_452), .CO(n_457), .S(n_456));
   FA_X1 i_229 (.A(n_454), .B(n_415), .CI(n_456), .CO(n_459), .S(n_458));
   HA_X1 i_230 (.A(n_417), .B(n_458), .CO(n_461), .S(n_460));
   FA_X1 i_231 (.A(p_0[23]), .B(p_1[23]), .CI(p_2[23]), .CO(n_463), .S(n_462));
   FA_X1 i_232 (.A(p_3[23]), .B(p_4[23]), .CI(p_5[23]), .CO(n_465), .S(n_464));
   FA_X1 i_233 (.A(p_6[23]), .B(p_7[23]), .CI(p_8[23]), .CO(n_467), .S(n_466));
   FA_X1 i_234 (.A(p_9[23]), .B(p_10[23]), .CI(p_11[23]), .CO(n_469), .S(n_468));
   FA_X1 i_235 (.A(p_12[23]), .B(p_13[23]), .CI(p_14[23]), .CO(n_471), .S(n_470));
   FA_X1 i_236 (.A(p_15[23]), .B(p_16[23]), .CI(p_17[23]), .CO(n_473), .S(n_472));
   FA_X1 i_237 (.A(p_18[23]), .B(p_19[23]), .CI(p_20[23]), .CO(n_475), .S(n_474));
   FA_X1 i_238 (.A(p_21[23]), .B(p_22[23]), .CI(out[23]), .CO(n_477), .S(n_476));
   FA_X1 i_239 (.A(n_433), .B(n_431), .CI(n_429), .CO(n_479), .S(n_478));
   FA_X1 i_240 (.A(n_427), .B(n_425), .CI(n_423), .CO(n_481), .S(n_480));
   FA_X1 i_241 (.A(n_421), .B(n_439), .CI(n_437), .CO(n_483), .S(n_482));
   FA_X1 i_242 (.A(n_435), .B(n_476), .CI(n_474), .CO(n_485), .S(n_484));
   FA_X1 i_243 (.A(n_472), .B(n_470), .CI(n_468), .CO(n_487), .S(n_486));
   FA_X1 i_244 (.A(n_466), .B(n_464), .CI(n_462), .CO(n_489), .S(n_488));
   FA_X1 i_245 (.A(n_480), .B(n_478), .CI(n_445), .CO(n_491), .S(n_490));
   FA_X1 i_246 (.A(n_443), .B(n_441), .CI(n_482), .CO(n_493), .S(n_492));
   FA_X1 i_247 (.A(n_449), .B(n_447), .CI(n_488), .CO(n_495), .S(n_494));
   FA_X1 i_248 (.A(n_486), .B(n_484), .CI(n_451), .CO(n_497), .S(n_496));
   FA_X1 i_249 (.A(n_492), .B(n_490), .CI(n_453), .CO(n_499), .S(n_498));
   FA_X1 i_250 (.A(n_494), .B(n_455), .CI(n_496), .CO(n_501), .S(n_500));
   FA_X1 i_251 (.A(n_498), .B(n_457), .CI(n_500), .CO(n_503), .S(n_502));
   HA_X1 i_252 (.A(n_459), .B(n_502), .CO(n_505), .S(n_504));
   FA_X1 i_253 (.A(p_0[24]), .B(p_1[24]), .CI(p_2[24]), .CO(n_507), .S(n_506));
   FA_X1 i_254 (.A(p_3[24]), .B(p_4[24]), .CI(p_5[24]), .CO(n_509), .S(n_508));
   FA_X1 i_255 (.A(p_6[24]), .B(p_7[24]), .CI(p_8[24]), .CO(n_511), .S(n_510));
   FA_X1 i_256 (.A(p_9[24]), .B(p_10[24]), .CI(p_11[24]), .CO(n_513), .S(n_512));
   FA_X1 i_257 (.A(p_12[24]), .B(p_13[24]), .CI(p_14[24]), .CO(n_515), .S(n_514));
   FA_X1 i_258 (.A(p_15[24]), .B(p_16[24]), .CI(p_17[24]), .CO(n_517), .S(n_516));
   FA_X1 i_259 (.A(p_18[24]), .B(p_19[24]), .CI(p_20[24]), .CO(n_519), .S(n_518));
   FA_X1 i_260 (.A(p_21[24]), .B(p_22[24]), .CI(p_23[24]), .CO(n_521), .S(n_520));
   FA_X1 i_261 (.A(out[24]), .B(n_477), .CI(n_475), .CO(n_523), .S(n_522));
   FA_X1 i_262 (.A(n_473), .B(n_471), .CI(n_469), .CO(n_525), .S(n_524));
   FA_X1 i_263 (.A(n_467), .B(n_465), .CI(n_463), .CO(n_527), .S(n_526));
   FA_X1 i_264 (.A(n_481), .B(n_479), .CI(n_520), .CO(n_529), .S(n_528));
   FA_X1 i_265 (.A(n_518), .B(n_516), .CI(n_514), .CO(n_531), .S(n_530));
   FA_X1 i_266 (.A(n_512), .B(n_510), .CI(n_508), .CO(n_533), .S(n_532));
   FA_X1 i_267 (.A(n_506), .B(n_483), .CI(n_526), .CO(n_535), .S(n_534));
   FA_X1 i_268 (.A(n_524), .B(n_522), .CI(n_489), .CO(n_537), .S(n_536));
   FA_X1 i_269 (.A(n_487), .B(n_485), .CI(n_528), .CO(n_539), .S(n_538));
   FA_X1 i_270 (.A(n_491), .B(n_532), .CI(n_530), .CO(n_541), .S(n_540));
   FA_X1 i_271 (.A(n_534), .B(n_493), .CI(n_538), .CO(n_543), .S(n_542));
   FA_X1 i_272 (.A(n_536), .B(n_495), .CI(n_497), .CO(n_545), .S(n_544));
   FA_X1 i_273 (.A(n_499), .B(n_540), .CI(n_542), .CO(n_547), .S(n_546));
   FA_X1 i_274 (.A(n_544), .B(n_501), .CI(n_546), .CO(n_549), .S(n_548));
   HA_X1 i_275 (.A(n_503), .B(n_548), .CO(n_551), .S(n_550));
   FA_X1 i_276 (.A(p_0[25]), .B(p_1[25]), .CI(p_2[25]), .CO(n_553), .S(n_552));
   FA_X1 i_277 (.A(p_3[25]), .B(p_4[25]), .CI(p_5[25]), .CO(n_555), .S(n_554));
   FA_X1 i_278 (.A(p_6[25]), .B(p_7[25]), .CI(p_8[25]), .CO(n_557), .S(n_556));
   FA_X1 i_279 (.A(p_9[25]), .B(p_10[25]), .CI(p_11[25]), .CO(n_559), .S(n_558));
   FA_X1 i_280 (.A(p_12[25]), .B(p_13[25]), .CI(p_14[25]), .CO(n_561), .S(n_560));
   FA_X1 i_281 (.A(p_15[25]), .B(p_16[25]), .CI(p_17[25]), .CO(n_563), .S(n_562));
   FA_X1 i_282 (.A(p_18[25]), .B(p_19[25]), .CI(p_20[25]), .CO(n_565), .S(n_564));
   FA_X1 i_283 (.A(p_21[25]), .B(p_22[25]), .CI(p_23[25]), .CO(n_567), .S(n_566));
   FA_X1 i_284 (.A(p_24[25]), .B(out[25]), .CI(n_521), .CO(n_569), .S(n_568));
   FA_X1 i_285 (.A(n_519), .B(n_517), .CI(n_515), .CO(n_571), .S(n_570));
   FA_X1 i_286 (.A(n_513), .B(n_511), .CI(n_509), .CO(n_573), .S(n_572));
   FA_X1 i_287 (.A(n_507), .B(n_527), .CI(n_525), .CO(n_575), .S(n_574));
   FA_X1 i_288 (.A(n_523), .B(n_568), .CI(n_566), .CO(n_577), .S(n_576));
   FA_X1 i_289 (.A(n_564), .B(n_562), .CI(n_560), .CO(n_579), .S(n_578));
   FA_X1 i_290 (.A(n_558), .B(n_556), .CI(n_554), .CO(n_581), .S(n_580));
   FA_X1 i_291 (.A(n_552), .B(n_572), .CI(n_570), .CO(n_583), .S(n_582));
   FA_X1 i_292 (.A(n_533), .B(n_531), .CI(n_529), .CO(n_585), .S(n_584));
   FA_X1 i_293 (.A(n_574), .B(n_537), .CI(n_535), .CO(n_587), .S(n_586));
   FA_X1 i_294 (.A(n_580), .B(n_578), .CI(n_576), .CO(n_589), .S(n_588));
   FA_X1 i_295 (.A(n_539), .B(n_584), .CI(n_582), .CO(n_591), .S(n_590));
   FA_X1 i_296 (.A(n_541), .B(n_586), .CI(n_543), .CO(n_593), .S(n_592));
   FA_X1 i_297 (.A(n_545), .B(n_588), .CI(n_590), .CO(n_595), .S(n_594));
   FA_X1 i_298 (.A(n_547), .B(n_592), .CI(n_594), .CO(n_597), .S(n_596));
   HA_X1 i_299 (.A(n_549), .B(n_551), .CO(n_599), .S(n_598));
   FA_X1 i_300 (.A(p_0[26]), .B(p_1[26]), .CI(p_2[26]), .CO(n_601), .S(n_600));
   FA_X1 i_301 (.A(p_3[26]), .B(p_4[26]), .CI(p_5[26]), .CO(n_603), .S(n_602));
   FA_X1 i_302 (.A(p_6[26]), .B(p_7[26]), .CI(p_8[26]), .CO(n_605), .S(n_604));
   FA_X1 i_303 (.A(p_9[26]), .B(p_10[26]), .CI(p_11[26]), .CO(n_607), .S(n_606));
   FA_X1 i_304 (.A(p_12[26]), .B(p_13[26]), .CI(p_14[26]), .CO(n_609), .S(n_608));
   FA_X1 i_305 (.A(p_15[26]), .B(p_16[26]), .CI(p_17[26]), .CO(n_611), .S(n_610));
   FA_X1 i_306 (.A(p_18[26]), .B(p_19[26]), .CI(p_20[26]), .CO(n_613), .S(n_612));
   FA_X1 i_307 (.A(p_21[26]), .B(p_22[26]), .CI(p_23[26]), .CO(n_615), .S(n_614));
   FA_X1 i_308 (.A(p_24[26]), .B(p_25[26]), .CI(out[26]), .CO(n_617), .S(n_616));
   FA_X1 i_309 (.A(n_567), .B(n_565), .CI(n_563), .CO(n_619), .S(n_618));
   FA_X1 i_310 (.A(n_561), .B(n_559), .CI(n_557), .CO(n_621), .S(n_620));
   FA_X1 i_311 (.A(n_555), .B(n_553), .CI(n_573), .CO(n_623), .S(n_622));
   FA_X1 i_312 (.A(n_571), .B(n_569), .CI(n_616), .CO(n_625), .S(n_624));
   FA_X1 i_313 (.A(n_614), .B(n_612), .CI(n_610), .CO(n_627), .S(n_626));
   FA_X1 i_314 (.A(n_608), .B(n_606), .CI(n_604), .CO(n_629), .S(n_628));
   FA_X1 i_315 (.A(n_602), .B(n_600), .CI(n_575), .CO(n_631), .S(n_630));
   FA_X1 i_316 (.A(n_622), .B(n_620), .CI(n_618), .CO(n_633), .S(n_632));
   FA_X1 i_317 (.A(n_581), .B(n_579), .CI(n_577), .CO(n_635), .S(n_634));
   FA_X1 i_318 (.A(n_624), .B(n_585), .CI(n_583), .CO(n_637), .S(n_636));
   FA_X1 i_319 (.A(n_630), .B(n_628), .CI(n_626), .CO(n_639), .S(n_638));
   FA_X1 i_320 (.A(n_587), .B(n_634), .CI(n_632), .CO(n_641), .S(n_640));
   FA_X1 i_321 (.A(n_589), .B(n_636), .CI(n_591), .CO(n_643), .S(n_642));
   FA_X1 i_322 (.A(n_638), .B(n_593), .CI(n_640), .CO(n_645), .S(n_644));
   FA_X1 i_323 (.A(n_642), .B(n_595), .CI(n_644), .CO(n_647), .S(n_646));
   HA_X1 i_324 (.A(n_597), .B(n_646), .CO(n_649), .S(n_648));
   FA_X1 i_325 (.A(p_0[27]), .B(p_1[27]), .CI(p_2[27]), .CO(n_651), .S(n_650));
   FA_X1 i_326 (.A(p_3[27]), .B(p_4[27]), .CI(p_5[27]), .CO(n_653), .S(n_652));
   FA_X1 i_327 (.A(p_6[27]), .B(p_7[27]), .CI(p_8[27]), .CO(n_655), .S(n_654));
   FA_X1 i_328 (.A(p_9[27]), .B(p_10[27]), .CI(p_11[27]), .CO(n_657), .S(n_656));
   FA_X1 i_329 (.A(p_12[27]), .B(p_13[27]), .CI(p_14[27]), .CO(n_659), .S(n_658));
   FA_X1 i_330 (.A(p_15[27]), .B(p_16[27]), .CI(p_17[27]), .CO(n_661), .S(n_660));
   FA_X1 i_331 (.A(p_18[27]), .B(p_19[27]), .CI(p_20[27]), .CO(n_663), .S(n_662));
   FA_X1 i_332 (.A(p_21[27]), .B(p_22[27]), .CI(p_23[27]), .CO(n_665), .S(n_664));
   FA_X1 i_333 (.A(p_24[27]), .B(p_25[27]), .CI(p_26[27]), .CO(n_667), .S(n_666));
   FA_X1 i_334 (.A(out[27]), .B(n_617), .CI(n_615), .CO(n_669), .S(n_668));
   FA_X1 i_335 (.A(n_613), .B(n_611), .CI(n_609), .CO(n_671), .S(n_670));
   FA_X1 i_336 (.A(n_607), .B(n_605), .CI(n_603), .CO(n_673), .S(n_672));
   FA_X1 i_337 (.A(n_601), .B(n_621), .CI(n_619), .CO(n_675), .S(n_674));
   FA_X1 i_338 (.A(n_666), .B(n_664), .CI(n_662), .CO(n_677), .S(n_676));
   FA_X1 i_339 (.A(n_660), .B(n_658), .CI(n_656), .CO(n_679), .S(n_678));
   FA_X1 i_340 (.A(n_654), .B(n_652), .CI(n_650), .CO(n_681), .S(n_680));
   FA_X1 i_341 (.A(n_623), .B(n_672), .CI(n_670), .CO(n_683), .S(n_682));
   FA_X1 i_342 (.A(n_668), .B(n_629), .CI(n_627), .CO(n_685), .S(n_684));
   FA_X1 i_343 (.A(n_625), .B(n_631), .CI(n_674), .CO(n_687), .S(n_686));
   FA_X1 i_344 (.A(n_635), .B(n_633), .CI(n_680), .CO(n_689), .S(n_688));
   FA_X1 i_345 (.A(n_678), .B(n_676), .CI(n_637), .CO(n_691), .S(n_690));
   FA_X1 i_346 (.A(n_684), .B(n_682), .CI(n_639), .CO(n_693), .S(n_692));
   FA_X1 i_347 (.A(n_686), .B(n_688), .CI(n_641), .CO(n_695), .S(n_694));
   FA_X1 i_348 (.A(n_690), .B(n_643), .CI(n_692), .CO(n_697), .S(n_696));
   FA_X1 i_349 (.A(n_694), .B(n_645), .CI(n_696), .CO(n_699), .S(n_698));
   HA_X1 i_350 (.A(n_647), .B(n_698), .CO(n_701), .S(n_700));
   FA_X1 i_351 (.A(p_0[28]), .B(p_1[28]), .CI(p_2[28]), .CO(n_703), .S(n_702));
   FA_X1 i_352 (.A(p_3[28]), .B(p_4[28]), .CI(p_5[28]), .CO(n_705), .S(n_704));
   FA_X1 i_353 (.A(p_6[28]), .B(p_7[28]), .CI(p_8[28]), .CO(n_707), .S(n_706));
   FA_X1 i_354 (.A(p_9[28]), .B(p_10[28]), .CI(p_11[28]), .CO(n_709), .S(n_708));
   FA_X1 i_355 (.A(p_12[28]), .B(p_13[28]), .CI(p_14[28]), .CO(n_711), .S(n_710));
   FA_X1 i_356 (.A(p_15[28]), .B(p_16[28]), .CI(p_17[28]), .CO(n_713), .S(n_712));
   FA_X1 i_357 (.A(p_18[28]), .B(p_19[28]), .CI(p_20[28]), .CO(n_715), .S(n_714));
   FA_X1 i_358 (.A(p_21[28]), .B(p_22[28]), .CI(p_23[28]), .CO(n_717), .S(n_716));
   FA_X1 i_359 (.A(p_24[28]), .B(p_25[28]), .CI(p_26[28]), .CO(n_719), .S(n_718));
   FA_X1 i_360 (.A(p_27[28]), .B(out[28]), .CI(n_667), .CO(n_721), .S(n_720));
   FA_X1 i_361 (.A(n_665), .B(n_663), .CI(n_661), .CO(n_723), .S(n_722));
   FA_X1 i_362 (.A(n_659), .B(n_657), .CI(n_655), .CO(n_725), .S(n_724));
   FA_X1 i_363 (.A(n_653), .B(n_651), .CI(n_673), .CO(n_727), .S(n_726));
   FA_X1 i_364 (.A(n_671), .B(n_669), .CI(n_720), .CO(n_729), .S(n_728));
   FA_X1 i_365 (.A(n_718), .B(n_716), .CI(n_714), .CO(n_731), .S(n_730));
   FA_X1 i_366 (.A(n_712), .B(n_710), .CI(n_708), .CO(n_733), .S(n_732));
   FA_X1 i_367 (.A(n_706), .B(n_704), .CI(n_702), .CO(n_735), .S(n_734));
   FA_X1 i_368 (.A(n_675), .B(n_726), .CI(n_724), .CO(n_737), .S(n_736));
   FA_X1 i_369 (.A(n_722), .B(n_681), .CI(n_679), .CO(n_739), .S(n_738));
   FA_X1 i_370 (.A(n_677), .B(n_728), .CI(n_685), .CO(n_741), .S(n_740));
   FA_X1 i_371 (.A(n_683), .B(n_734), .CI(n_732), .CO(n_743), .S(n_742));
   FA_X1 i_372 (.A(n_730), .B(n_687), .CI(n_738), .CO(n_745), .S(n_744));
   FA_X1 i_373 (.A(n_736), .B(n_689), .CI(n_691), .CO(n_747), .S(n_746));
   FA_X1 i_374 (.A(n_740), .B(n_693), .CI(n_742), .CO(n_749), .S(n_748));
   FA_X1 i_375 (.A(n_744), .B(n_695), .CI(n_746), .CO(n_751), .S(n_750));
   FA_X1 i_376 (.A(n_748), .B(n_697), .CI(n_750), .CO(n_753), .S(n_752));
   HA_X1 i_377 (.A(n_699), .B(n_752), .CO(n_755), .S(n_754));
   FA_X1 i_378 (.A(p_0[29]), .B(p_1[29]), .CI(p_2[29]), .CO(n_757), .S(n_756));
   FA_X1 i_379 (.A(p_3[29]), .B(p_4[29]), .CI(p_5[29]), .CO(n_759), .S(n_758));
   FA_X1 i_380 (.A(p_6[29]), .B(p_7[29]), .CI(p_8[29]), .CO(n_761), .S(n_760));
   FA_X1 i_381 (.A(p_9[29]), .B(p_10[29]), .CI(p_11[29]), .CO(n_763), .S(n_762));
   FA_X1 i_382 (.A(p_12[29]), .B(p_13[29]), .CI(p_14[29]), .CO(n_765), .S(n_764));
   FA_X1 i_383 (.A(p_15[29]), .B(p_16[29]), .CI(p_17[29]), .CO(n_767), .S(n_766));
   FA_X1 i_384 (.A(p_18[29]), .B(p_19[29]), .CI(p_20[29]), .CO(n_769), .S(n_768));
   FA_X1 i_385 (.A(p_21[29]), .B(p_22[29]), .CI(p_23[29]), .CO(n_771), .S(n_770));
   FA_X1 i_386 (.A(p_24[29]), .B(p_25[29]), .CI(p_26[29]), .CO(n_773), .S(n_772));
   FA_X1 i_387 (.A(p_27[29]), .B(p_28[29]), .CI(out[29]), .CO(n_775), .S(n_774));
   FA_X1 i_388 (.A(n_719), .B(n_717), .CI(n_715), .CO(n_777), .S(n_776));
   FA_X1 i_389 (.A(n_713), .B(n_711), .CI(n_709), .CO(n_779), .S(n_778));
   FA_X1 i_390 (.A(n_707), .B(n_705), .CI(n_703), .CO(n_781), .S(n_780));
   FA_X1 i_391 (.A(n_725), .B(n_723), .CI(n_721), .CO(n_783), .S(n_782));
   FA_X1 i_392 (.A(n_774), .B(n_772), .CI(n_770), .CO(n_785), .S(n_784));
   FA_X1 i_393 (.A(n_768), .B(n_766), .CI(n_764), .CO(n_787), .S(n_786));
   FA_X1 i_394 (.A(n_762), .B(n_760), .CI(n_758), .CO(n_789), .S(n_788));
   FA_X1 i_395 (.A(n_756), .B(n_727), .CI(n_780), .CO(n_791), .S(n_790));
   FA_X1 i_396 (.A(n_778), .B(n_776), .CI(n_735), .CO(n_793), .S(n_792));
   FA_X1 i_397 (.A(n_733), .B(n_731), .CI(n_729), .CO(n_795), .S(n_794));
   FA_X1 i_398 (.A(n_782), .B(n_739), .CI(n_737), .CO(n_797), .S(n_796));
   FA_X1 i_399 (.A(n_788), .B(n_786), .CI(n_784), .CO(n_799), .S(n_798));
   FA_X1 i_400 (.A(n_790), .B(n_741), .CI(n_794), .CO(n_801), .S(n_800));
   FA_X1 i_401 (.A(n_792), .B(n_743), .CI(n_796), .CO(n_803), .S(n_802));
   FA_X1 i_402 (.A(n_745), .B(n_747), .CI(n_798), .CO(n_805), .S(n_804));
   FA_X1 i_403 (.A(n_800), .B(n_802), .CI(n_749), .CO(n_807), .S(n_806));
   FA_X1 i_404 (.A(n_751), .B(n_804), .CI(n_806), .CO(n_809), .S(n_808));
   HA_X1 i_405 (.A(n_753), .B(n_808), .CO(n_811), .S(n_810));
   FA_X1 i_406 (.A(p_0[30]), .B(p_1[30]), .CI(p_2[30]), .CO(n_813), .S(n_812));
   FA_X1 i_407 (.A(p_3[30]), .B(p_4[30]), .CI(p_5[30]), .CO(n_815), .S(n_814));
   FA_X1 i_408 (.A(p_6[30]), .B(p_7[30]), .CI(p_8[30]), .CO(n_817), .S(n_816));
   FA_X1 i_409 (.A(p_9[30]), .B(p_10[30]), .CI(p_11[30]), .CO(n_819), .S(n_818));
   FA_X1 i_410 (.A(p_12[30]), .B(p_13[30]), .CI(p_14[30]), .CO(n_821), .S(n_820));
   FA_X1 i_411 (.A(p_15[30]), .B(p_16[30]), .CI(p_17[30]), .CO(n_823), .S(n_822));
   FA_X1 i_412 (.A(p_18[30]), .B(p_19[30]), .CI(p_20[30]), .CO(n_825), .S(n_824));
   FA_X1 i_413 (.A(p_21[30]), .B(p_22[30]), .CI(p_23[30]), .CO(n_827), .S(n_826));
   FA_X1 i_414 (.A(p_24[30]), .B(p_25[30]), .CI(p_26[30]), .CO(n_829), .S(n_828));
   FA_X1 i_415 (.A(p_27[30]), .B(p_28[30]), .CI(p_29[30]), .CO(n_831), .S(n_830));
   FA_X1 i_416 (.A(out[30]), .B(n_775), .CI(n_773), .CO(n_833), .S(n_832));
   FA_X1 i_417 (.A(n_771), .B(n_769), .CI(n_767), .CO(n_835), .S(n_834));
   FA_X1 i_418 (.A(n_765), .B(n_763), .CI(n_761), .CO(n_837), .S(n_836));
   FA_X1 i_419 (.A(n_759), .B(n_757), .CI(n_781), .CO(n_839), .S(n_838));
   FA_X1 i_420 (.A(n_779), .B(n_777), .CI(n_830), .CO(n_841), .S(n_840));
   FA_X1 i_421 (.A(n_828), .B(n_826), .CI(n_824), .CO(n_843), .S(n_842));
   FA_X1 i_422 (.A(n_822), .B(n_820), .CI(n_818), .CO(n_845), .S(n_844));
   FA_X1 i_423 (.A(n_816), .B(n_814), .CI(n_812), .CO(n_847), .S(n_846));
   FA_X1 i_424 (.A(n_783), .B(n_838), .CI(n_836), .CO(n_849), .S(n_848));
   FA_X1 i_425 (.A(n_834), .B(n_832), .CI(n_789), .CO(n_851), .S(n_850));
   FA_X1 i_426 (.A(n_787), .B(n_785), .CI(n_840), .CO(n_853), .S(n_852));
   FA_X1 i_427 (.A(n_795), .B(n_793), .CI(n_791), .CO(n_855), .S(n_854));
   FA_X1 i_428 (.A(n_846), .B(n_844), .CI(n_842), .CO(n_857), .S(n_856));
   FA_X1 i_429 (.A(n_797), .B(n_852), .CI(n_850), .CO(n_859), .S(n_858));
   FA_X1 i_430 (.A(n_848), .B(n_799), .CI(n_854), .CO(n_861), .S(n_860));
   FA_X1 i_431 (.A(n_801), .B(n_856), .CI(n_803), .CO(n_863), .S(n_862));
   FA_X1 i_432 (.A(n_860), .B(n_858), .CI(n_805), .CO(n_865), .S(n_864));
   FA_X1 i_433 (.A(n_807), .B(n_862), .CI(n_864), .CO(n_867), .S(n_866));
   HA_X1 i_434 (.A(n_809), .B(n_866), .CO(n_869), .S(n_868));
   FA_X1 i_435 (.A(p_0[31]), .B(p_1[31]), .CI(p_2[31]), .CO(n_871), .S(n_870));
   FA_X1 i_436 (.A(p_3[31]), .B(p_4[31]), .CI(p_5[31]), .CO(n_873), .S(n_872));
   FA_X1 i_437 (.A(p_6[31]), .B(p_7[31]), .CI(p_8[31]), .CO(n_875), .S(n_874));
   FA_X1 i_438 (.A(p_9[31]), .B(p_10[31]), .CI(p_11[31]), .CO(n_877), .S(n_876));
   FA_X1 i_439 (.A(p_12[31]), .B(p_13[31]), .CI(p_14[31]), .CO(n_879), .S(n_878));
   FA_X1 i_440 (.A(p_15[31]), .B(p_16[31]), .CI(p_17[31]), .CO(n_881), .S(n_880));
   FA_X1 i_441 (.A(p_18[31]), .B(p_19[31]), .CI(p_20[31]), .CO(n_883), .S(n_882));
   FA_X1 i_442 (.A(p_21[31]), .B(p_22[31]), .CI(p_23[31]), .CO(n_885), .S(n_884));
   FA_X1 i_443 (.A(p_24[31]), .B(p_25[31]), .CI(p_26[31]), .CO(n_887), .S(n_886));
   FA_X1 i_444 (.A(p_27[31]), .B(p_28[31]), .CI(p_29[31]), .CO(n_889), .S(n_888));
   FA_X1 i_445 (.A(p_30[31]), .B(out[31]), .CI(n_831), .CO(n_891), .S(n_890));
   FA_X1 i_446 (.A(n_829), .B(n_827), .CI(n_825), .CO(n_893), .S(n_892));
   FA_X1 i_447 (.A(n_823), .B(n_821), .CI(n_819), .CO(n_895), .S(n_894));
   FA_X1 i_448 (.A(n_817), .B(n_815), .CI(n_813), .CO(n_897), .S(n_896));
   FA_X1 i_449 (.A(n_837), .B(n_835), .CI(n_833), .CO(n_899), .S(n_898));
   FA_X1 i_450 (.A(n_890), .B(n_888), .CI(n_886), .CO(n_901), .S(n_900));
   FA_X1 i_451 (.A(n_884), .B(n_882), .CI(n_880), .CO(n_903), .S(n_902));
   FA_X1 i_452 (.A(n_878), .B(n_876), .CI(n_874), .CO(n_905), .S(n_904));
   FA_X1 i_453 (.A(n_872), .B(n_870), .CI(n_839), .CO(n_907), .S(n_906));
   FA_X1 i_454 (.A(n_896), .B(n_894), .CI(n_892), .CO(n_909), .S(n_908));
   FA_X1 i_455 (.A(n_847), .B(n_845), .CI(n_843), .CO(n_911), .S(n_910));
   FA_X1 i_456 (.A(n_841), .B(n_898), .CI(n_851), .CO(n_913), .S(n_912));
   FA_X1 i_457 (.A(n_849), .B(n_906), .CI(n_904), .CO(n_915), .S(n_914));
   FA_X1 i_458 (.A(n_902), .B(n_900), .CI(n_855), .CO(n_917), .S(n_916));
   FA_X1 i_459 (.A(n_853), .B(n_910), .CI(n_908), .CO(n_919), .S(n_918));
   FA_X1 i_460 (.A(n_857), .B(n_912), .CI(n_859), .CO(n_921), .S(n_920));
   FA_X1 i_461 (.A(n_916), .B(n_914), .CI(n_861), .CO(n_923), .S(n_922));
   FA_X1 i_462 (.A(n_918), .B(n_863), .CI(n_920), .CO(n_925), .S(n_924));
   FA_X1 i_463 (.A(n_865), .B(n_922), .CI(n_924), .CO(n_927), .S(n_926));
   HA_X1 i_464 (.A(n_867), .B(n_926), .CO(n_929), .S(n_928));
   FA_X1 i_465 (.A(p_2[32]), .B(p_3[32]), .CI(p_4[32]), .CO(n_931), .S(n_930));
   FA_X1 i_466 (.A(p_5[32]), .B(p_6[32]), .CI(p_7[32]), .CO(n_933), .S(n_932));
   FA_X1 i_467 (.A(p_8[32]), .B(p_9[32]), .CI(p_10[32]), .CO(n_935), .S(n_934));
   FA_X1 i_468 (.A(p_11[32]), .B(p_12[32]), .CI(p_13[32]), .CO(n_937), .S(n_936));
   FA_X1 i_469 (.A(p_14[32]), .B(p_15[32]), .CI(p_16[32]), .CO(n_939), .S(n_938));
   FA_X1 i_470 (.A(p_17[32]), .B(p_18[32]), .CI(p_19[32]), .CO(n_941), .S(n_940));
   FA_X1 i_471 (.A(p_20[32]), .B(p_21[32]), .CI(p_22[32]), .CO(n_943), .S(n_942));
   FA_X1 i_472 (.A(p_23[32]), .B(p_24[32]), .CI(p_25[32]), .CO(n_945), .S(n_944));
   FA_X1 i_473 (.A(p_26[32]), .B(p_27[32]), .CI(p_28[32]), .CO(n_947), .S(n_946));
   FA_X1 i_474 (.A(n_889), .B(n_887), .CI(n_885), .CO(n_949), .S(n_948));
   FA_X1 i_475 (.A(n_883), .B(n_881), .CI(n_879), .CO(n_951), .S(n_950));
   FA_X1 i_476 (.A(n_877), .B(n_875), .CI(n_873), .CO(n_953), .S(n_952));
   FA_X1 i_477 (.A(n_871), .B(n_897), .CI(n_895), .CO(n_955), .S(n_954));
   FA_X1 i_478 (.A(n_893), .B(n_891), .CI(n_1944), .CO(n_957), .S(n_956));
   FA_X1 i_479 (.A(n_946), .B(n_944), .CI(n_942), .CO(n_959), .S(n_958));
   FA_X1 i_480 (.A(n_940), .B(n_938), .CI(n_936), .CO(n_961), .S(n_960));
   FA_X1 i_481 (.A(n_934), .B(n_932), .CI(n_930), .CO(n_963), .S(n_962));
   FA_X1 i_482 (.A(n_1949), .B(n_899), .CI(n_952), .CO(n_965), .S(n_964));
   FA_X1 i_483 (.A(n_950), .B(n_948), .CI(n_905), .CO(n_967), .S(n_966));
   FA_X1 i_484 (.A(n_903), .B(n_901), .CI(n_907), .CO(n_969), .S(n_968));
   FA_X1 i_485 (.A(n_956), .B(n_954), .CI(n_911), .CO(n_971), .S(n_970));
   FA_X1 i_486 (.A(n_909), .B(n_962), .CI(n_960), .CO(n_973), .S(n_972));
   FA_X1 i_487 (.A(n_958), .B(n_964), .CI(n_913), .CO(n_975), .S(n_974));
   FA_X1 i_488 (.A(n_968), .B(n_966), .CI(n_915), .CO(n_977), .S(n_976));
   FA_X1 i_489 (.A(n_917), .B(n_970), .CI(n_919), .CO(n_979), .S(n_978));
   FA_X1 i_490 (.A(n_972), .B(n_974), .CI(n_921), .CO(n_981), .S(n_980));
   FA_X1 i_491 (.A(n_976), .B(n_923), .CI(n_978), .CO(n_983), .S(n_982));
   FA_X1 i_492 (.A(n_980), .B(n_925), .CI(n_982), .CO(n_985), .S(n_984));
   HA_X1 i_493 (.A(n_927), .B(n_984), .CO(n_987), .S(n_986));
   FA_X1 i_494 (.A(p_3[33]), .B(p_4[33]), .CI(p_5[33]), .CO(n_989), .S(n_988));
   FA_X1 i_495 (.A(p_6[33]), .B(p_7[33]), .CI(p_8[33]), .CO(n_991), .S(n_990));
   FA_X1 i_496 (.A(p_9[33]), .B(p_10[33]), .CI(p_11[33]), .CO(n_993), .S(n_992));
   FA_X1 i_497 (.A(p_12[33]), .B(p_13[33]), .CI(p_14[33]), .CO(n_995), .S(n_994));
   FA_X1 i_498 (.A(p_15[33]), .B(p_16[33]), .CI(p_17[33]), .CO(n_997), .S(n_996));
   FA_X1 i_499 (.A(p_18[33]), .B(p_19[33]), .CI(p_20[33]), .CO(n_999), .S(n_998));
   FA_X1 i_500 (.A(p_21[33]), .B(p_22[33]), .CI(p_23[33]), .CO(n_1001), .S(
      n_1000));
   FA_X1 i_501 (.A(p_24[33]), .B(p_25[33]), .CI(p_26[33]), .CO(n_1003), .S(
      n_1002));
   FA_X1 i_502 (.A(p_27[33]), .B(p_28[33]), .CI(p_29[33]), .CO(n_1005), .S(
      n_1004));
   FA_X1 i_503 (.A(p_30[33]), .B(n_1946), .CI(n_947), .CO(n_1007), .S(n_1006));
   FA_X1 i_504 (.A(n_945), .B(n_943), .CI(n_941), .CO(n_1009), .S(n_1008));
   FA_X1 i_505 (.A(n_939), .B(n_937), .CI(n_935), .CO(n_1011), .S(n_1010));
   FA_X1 i_506 (.A(n_933), .B(n_931), .CI(n_1950), .CO(n_1013), .S(n_1012));
   FA_X1 i_507 (.A(n_953), .B(n_951), .CI(n_949), .CO(n_1015), .S(n_1014));
   FA_X1 i_508 (.A(n_1004), .B(n_1002), .CI(n_1000), .CO(n_1017), .S(n_1016));
   FA_X1 i_509 (.A(n_998), .B(n_996), .CI(n_994), .CO(n_1019), .S(n_1018));
   FA_X1 i_510 (.A(n_992), .B(n_990), .CI(n_988), .CO(n_1021), .S(n_1020));
   FA_X1 i_511 (.A(n_1941), .B(n_955), .CI(n_1012), .CO(n_1023), .S(n_1022));
   FA_X1 i_512 (.A(n_1010), .B(n_1008), .CI(n_1006), .CO(n_1025), .S(n_1024));
   FA_X1 i_513 (.A(n_963), .B(n_961), .CI(n_959), .CO(n_1027), .S(n_1026));
   FA_X1 i_514 (.A(n_957), .B(n_1014), .CI(n_967), .CO(n_1029), .S(n_1028));
   FA_X1 i_515 (.A(n_965), .B(n_969), .CI(n_1020), .CO(n_1031), .S(n_1030));
   FA_X1 i_516 (.A(n_1018), .B(n_1016), .CI(n_1022), .CO(n_1033), .S(n_1032));
   FA_X1 i_517 (.A(n_971), .B(n_1026), .CI(n_1024), .CO(n_1035), .S(n_1034));
   FA_X1 i_518 (.A(n_973), .B(n_975), .CI(n_1028), .CO(n_1037), .S(n_1036));
   FA_X1 i_519 (.A(n_977), .B(n_1030), .CI(n_1032), .CO(n_1039), .S(n_1038));
   FA_X1 i_520 (.A(n_979), .B(n_1034), .CI(n_1036), .CO(n_1041), .S(n_1040));
   FA_X1 i_521 (.A(n_981), .B(n_1038), .CI(n_983), .CO(n_1043), .S(n_1042));
   FA_X1 i_522 (.A(n_1040), .B(n_1042), .CI(n_985), .CO(n_1045), .S(n_1044));
   FA_X1 i_523 (.A(p_4[34]), .B(p_5[34]), .CI(p_6[34]), .CO(n_1047), .S(n_1046));
   FA_X1 i_524 (.A(p_7[34]), .B(p_8[34]), .CI(p_9[34]), .CO(n_1049), .S(n_1048));
   FA_X1 i_525 (.A(p_10[34]), .B(p_11[34]), .CI(p_12[34]), .CO(n_1051), .S(
      n_1050));
   FA_X1 i_526 (.A(p_13[34]), .B(p_14[34]), .CI(p_15[34]), .CO(n_1053), .S(
      n_1052));
   FA_X1 i_527 (.A(p_16[34]), .B(p_17[34]), .CI(p_18[34]), .CO(n_1055), .S(
      n_1054));
   FA_X1 i_528 (.A(p_19[34]), .B(p_20[34]), .CI(p_21[34]), .CO(n_1057), .S(
      n_1056));
   FA_X1 i_529 (.A(p_22[34]), .B(p_23[34]), .CI(p_24[34]), .CO(n_1059), .S(
      n_1058));
   FA_X1 i_530 (.A(p_25[34]), .B(p_26[34]), .CI(p_27[34]), .CO(n_1061), .S(
      n_1060));
   FA_X1 i_531 (.A(p_28[34]), .B(p_29[34]), .CI(p_30[34]), .CO(n_1063), .S(
      n_1062));
   FA_X1 i_532 (.A(n_1005), .B(n_1003), .CI(n_1001), .CO(n_1065), .S(n_1064));
   FA_X1 i_533 (.A(n_999), .B(n_997), .CI(n_995), .CO(n_1067), .S(n_1066));
   FA_X1 i_534 (.A(n_993), .B(n_991), .CI(n_989), .CO(n_1069), .S(n_1068));
   FA_X1 i_535 (.A(n_1943), .B(n_1013), .CI(n_1011), .CO(n_1071), .S(n_1070));
   FA_X1 i_536 (.A(n_1009), .B(n_1007), .CI(n_1062), .CO(n_1073), .S(n_1072));
   FA_X1 i_537 (.A(n_1060), .B(n_1058), .CI(n_1056), .CO(n_1075), .S(n_1074));
   FA_X1 i_538 (.A(n_1054), .B(n_1052), .CI(n_1050), .CO(n_1077), .S(n_1076));
   FA_X1 i_539 (.A(n_1048), .B(n_1046), .CI(n_1938), .CO(n_1079), .S(n_1078));
   FA_X1 i_540 (.A(n_1015), .B(n_1068), .CI(n_1066), .CO(n_1081), .S(n_1080));
   FA_X1 i_541 (.A(n_1064), .B(n_1021), .CI(n_1019), .CO(n_1083), .S(n_1082));
   FA_X1 i_542 (.A(n_1017), .B(n_1072), .CI(n_1070), .CO(n_1085), .S(n_1084));
   FA_X1 i_543 (.A(n_1027), .B(n_1025), .CI(n_1023), .CO(n_1087), .S(n_1086));
   FA_X1 i_544 (.A(n_1078), .B(n_1076), .CI(n_1074), .CO(n_1089), .S(n_1088));
   FA_X1 i_545 (.A(n_1029), .B(n_1082), .CI(n_1080), .CO(n_1091), .S(n_1090));
   FA_X1 i_546 (.A(n_1031), .B(n_1033), .CI(n_1086), .CO(n_1093), .S(n_1092));
   FA_X1 i_547 (.A(n_1084), .B(n_1035), .CI(n_1088), .CO(n_1095), .S(n_1094));
   FA_X1 i_548 (.A(n_1037), .B(n_1090), .CI(n_1039), .CO(n_1097), .S(n_1096));
   FA_X1 i_549 (.A(n_1092), .B(n_1094), .CI(n_1041), .CO(n_1099), .S(n_1098));
   FA_X1 i_550 (.A(n_1096), .B(n_1043), .CI(n_1098), .CO(n_1101), .S(n_1100));
   FA_X1 i_551 (.A(p_5[35]), .B(p_6[35]), .CI(p_7[35]), .CO(n_1103), .S(n_1102));
   FA_X1 i_552 (.A(p_8[35]), .B(p_9[35]), .CI(p_10[35]), .CO(n_1105), .S(n_1104));
   FA_X1 i_553 (.A(p_11[35]), .B(p_12[35]), .CI(p_13[35]), .CO(n_1107), .S(
      n_1106));
   FA_X1 i_554 (.A(p_14[35]), .B(p_15[35]), .CI(p_16[35]), .CO(n_1109), .S(
      n_1108));
   FA_X1 i_555 (.A(p_17[35]), .B(p_18[35]), .CI(p_19[35]), .CO(n_1111), .S(
      n_1110));
   FA_X1 i_556 (.A(p_20[35]), .B(p_21[35]), .CI(p_22[35]), .CO(n_1113), .S(
      n_1112));
   FA_X1 i_557 (.A(p_23[35]), .B(p_24[35]), .CI(p_25[35]), .CO(n_1115), .S(
      n_1114));
   FA_X1 i_558 (.A(p_26[35]), .B(p_27[35]), .CI(p_28[35]), .CO(n_1117), .S(
      n_1116));
   FA_X1 i_559 (.A(p_29[35]), .B(p_30[35]), .CI(n_1063), .CO(n_1119), .S(n_1118));
   FA_X1 i_560 (.A(n_1061), .B(n_1059), .CI(n_1057), .CO(n_1121), .S(n_1120));
   FA_X1 i_561 (.A(n_1055), .B(n_1053), .CI(n_1051), .CO(n_1123), .S(n_1122));
   FA_X1 i_562 (.A(n_1049), .B(n_1047), .CI(n_1940), .CO(n_1125), .S(n_1124));
   FA_X1 i_563 (.A(n_1069), .B(n_1067), .CI(n_1065), .CO(n_1127), .S(n_1126));
   FA_X1 i_564 (.A(n_1118), .B(n_1116), .CI(n_1114), .CO(n_1129), .S(n_1128));
   FA_X1 i_565 (.A(n_1112), .B(n_1110), .CI(n_1108), .CO(n_1131), .S(n_1130));
   FA_X1 i_566 (.A(n_1106), .B(n_1104), .CI(n_1102), .CO(n_1133), .S(n_1132));
   FA_X1 i_567 (.A(n_1935), .B(n_1071), .CI(n_1124), .CO(n_1135), .S(n_1134));
   FA_X1 i_568 (.A(n_1122), .B(n_1120), .CI(n_1079), .CO(n_1137), .S(n_1136));
   FA_X1 i_569 (.A(n_1077), .B(n_1075), .CI(n_1073), .CO(n_1139), .S(n_1138));
   FA_X1 i_570 (.A(n_1126), .B(n_1083), .CI(n_1081), .CO(n_1141), .S(n_1140));
   FA_X1 i_571 (.A(n_1132), .B(n_1130), .CI(n_1128), .CO(n_1143), .S(n_1142));
   FA_X1 i_572 (.A(n_1134), .B(n_1087), .CI(n_1085), .CO(n_1145), .S(n_1144));
   FA_X1 i_573 (.A(n_1138), .B(n_1136), .CI(n_1089), .CO(n_1147), .S(n_1146));
   FA_X1 i_574 (.A(n_1140), .B(n_1091), .CI(n_1142), .CO(n_1149), .S(n_1148));
   FA_X1 i_575 (.A(n_1144), .B(n_1093), .CI(n_1146), .CO(n_1151), .S(n_1150));
   FA_X1 i_576 (.A(n_1095), .B(n_1148), .CI(n_1097), .CO(n_1153), .S(n_1152));
   FA_X1 i_577 (.A(n_1150), .B(n_1099), .CI(n_1152), .CO(n_1155), .S(n_1154));
   FA_X1 i_578 (.A(p_6[36]), .B(p_7[36]), .CI(p_8[36]), .CO(n_1157), .S(n_1156));
   FA_X1 i_579 (.A(p_9[36]), .B(p_10[36]), .CI(p_11[36]), .CO(n_1159), .S(n_1158));
   FA_X1 i_580 (.A(p_12[36]), .B(p_13[36]), .CI(p_14[36]), .CO(n_1161), .S(
      n_1160));
   FA_X1 i_581 (.A(p_15[36]), .B(p_16[36]), .CI(p_17[36]), .CO(n_1163), .S(
      n_1162));
   FA_X1 i_582 (.A(p_18[36]), .B(p_19[36]), .CI(p_20[36]), .CO(n_1165), .S(
      n_1164));
   FA_X1 i_583 (.A(p_21[36]), .B(p_22[36]), .CI(p_23[36]), .CO(n_1167), .S(
      n_1166));
   FA_X1 i_584 (.A(p_24[36]), .B(p_25[36]), .CI(p_26[36]), .CO(n_1169), .S(
      n_1168));
   FA_X1 i_585 (.A(p_27[36]), .B(p_28[36]), .CI(p_29[36]), .CO(n_1171), .S(
      n_1170));
   FA_X1 i_586 (.A(p_30[36]), .B(n_1117), .CI(n_1115), .CO(n_1173), .S(n_1172));
   FA_X1 i_587 (.A(n_1113), .B(n_1111), .CI(n_1109), .CO(n_1175), .S(n_1174));
   FA_X1 i_588 (.A(n_1107), .B(n_1105), .CI(n_1103), .CO(n_1177), .S(n_1176));
   FA_X1 i_589 (.A(n_1937), .B(n_1125), .CI(n_1123), .CO(n_1179), .S(n_1178));
   FA_X1 i_590 (.A(n_1121), .B(n_1119), .CI(n_1170), .CO(n_1181), .S(n_1180));
   FA_X1 i_591 (.A(n_1168), .B(n_1166), .CI(n_1164), .CO(n_1183), .S(n_1182));
   FA_X1 i_592 (.A(n_1162), .B(n_1160), .CI(n_1158), .CO(n_1185), .S(n_1184));
   FA_X1 i_593 (.A(n_1156), .B(n_1932), .CI(n_1127), .CO(n_1187), .S(n_1186));
   FA_X1 i_594 (.A(n_1176), .B(n_1174), .CI(n_1172), .CO(n_1189), .S(n_1188));
   FA_X1 i_595 (.A(n_1133), .B(n_1131), .CI(n_1129), .CO(n_1191), .S(n_1190));
   FA_X1 i_596 (.A(n_1180), .B(n_1178), .CI(n_1139), .CO(n_1193), .S(n_1192));
   FA_X1 i_597 (.A(n_1137), .B(n_1135), .CI(n_1186), .CO(n_1195), .S(n_1194));
   FA_X1 i_598 (.A(n_1184), .B(n_1182), .CI(n_1141), .CO(n_1197), .S(n_1196));
   FA_X1 i_599 (.A(n_1190), .B(n_1188), .CI(n_1143), .CO(n_1199), .S(n_1198));
   FA_X1 i_600 (.A(n_1145), .B(n_1194), .CI(n_1192), .CO(n_1201), .S(n_1200));
   FA_X1 i_601 (.A(n_1147), .B(n_1196), .CI(n_1198), .CO(n_1203), .S(n_1202));
   FA_X1 i_602 (.A(n_1149), .B(n_1200), .CI(n_1151), .CO(n_1205), .S(n_1204));
   FA_X1 i_603 (.A(n_1202), .B(n_1153), .CI(n_1204), .CO(n_1207), .S(n_1206));
   FA_X1 i_604 (.A(p_7[37]), .B(p_8[37]), .CI(p_9[37]), .CO(n_1209), .S(n_1208));
   FA_X1 i_605 (.A(p_10[37]), .B(p_11[37]), .CI(p_12[37]), .CO(n_1211), .S(
      n_1210));
   FA_X1 i_606 (.A(p_13[37]), .B(p_14[37]), .CI(p_15[37]), .CO(n_1213), .S(
      n_1212));
   FA_X1 i_607 (.A(p_16[37]), .B(p_17[37]), .CI(p_18[37]), .CO(n_1215), .S(
      n_1214));
   FA_X1 i_608 (.A(p_19[37]), .B(p_20[37]), .CI(p_21[37]), .CO(n_1217), .S(
      n_1216));
   FA_X1 i_609 (.A(p_22[37]), .B(p_23[37]), .CI(p_24[37]), .CO(n_1219), .S(
      n_1218));
   FA_X1 i_610 (.A(p_25[37]), .B(p_26[37]), .CI(p_27[37]), .CO(n_1221), .S(
      n_1220));
   FA_X1 i_611 (.A(p_28[37]), .B(p_29[37]), .CI(p_30[37]), .CO(n_1223), .S(
      n_1222));
   FA_X1 i_612 (.A(n_1171), .B(n_1169), .CI(n_1167), .CO(n_1225), .S(n_1224));
   FA_X1 i_613 (.A(n_1165), .B(n_1163), .CI(n_1161), .CO(n_1227), .S(n_1226));
   FA_X1 i_614 (.A(n_1159), .B(n_1157), .CI(n_1934), .CO(n_1229), .S(n_1228));
   FA_X1 i_615 (.A(n_1177), .B(n_1175), .CI(n_1173), .CO(n_1231), .S(n_1230));
   FA_X1 i_616 (.A(n_1222), .B(n_1220), .CI(n_1218), .CO(n_1233), .S(n_1232));
   FA_X1 i_617 (.A(n_1216), .B(n_1214), .CI(n_1212), .CO(n_1235), .S(n_1234));
   FA_X1 i_618 (.A(n_1210), .B(n_1208), .CI(n_1929), .CO(n_1237), .S(n_1236));
   FA_X1 i_619 (.A(n_1179), .B(n_1228), .CI(n_1226), .CO(n_1239), .S(n_1238));
   FA_X1 i_620 (.A(n_1224), .B(n_1185), .CI(n_1183), .CO(n_1241), .S(n_1240));
   FA_X1 i_621 (.A(n_1181), .B(n_1187), .CI(n_1230), .CO(n_1243), .S(n_1242));
   FA_X1 i_622 (.A(n_1191), .B(n_1189), .CI(n_1236), .CO(n_1245), .S(n_1244));
   FA_X1 i_623 (.A(n_1234), .B(n_1232), .CI(n_1193), .CO(n_1247), .S(n_1246));
   FA_X1 i_624 (.A(n_1240), .B(n_1238), .CI(n_1195), .CO(n_1249), .S(n_1248));
   FA_X1 i_625 (.A(n_1242), .B(n_1197), .CI(n_1244), .CO(n_1251), .S(n_1250));
   FA_X1 i_626 (.A(n_1199), .B(n_1246), .CI(n_1201), .CO(n_1253), .S(n_1252));
   FA_X1 i_627 (.A(n_1248), .B(n_1250), .CI(n_1203), .CO(n_1255), .S(n_1254));
   FA_X1 i_628 (.A(n_1252), .B(n_1205), .CI(n_1254), .CO(n_1257), .S(n_1256));
   FA_X1 i_629 (.A(p_8[38]), .B(p_9[38]), .CI(p_10[38]), .CO(n_1259), .S(n_1258));
   FA_X1 i_630 (.A(p_11[38]), .B(p_12[38]), .CI(p_13[38]), .CO(n_1261), .S(
      n_1260));
   FA_X1 i_631 (.A(p_14[38]), .B(p_15[38]), .CI(p_16[38]), .CO(n_1263), .S(
      n_1262));
   FA_X1 i_632 (.A(p_17[38]), .B(p_18[38]), .CI(p_19[38]), .CO(n_1265), .S(
      n_1264));
   FA_X1 i_633 (.A(p_20[38]), .B(p_21[38]), .CI(p_22[38]), .CO(n_1267), .S(
      n_1266));
   FA_X1 i_634 (.A(p_23[38]), .B(p_24[38]), .CI(p_25[38]), .CO(n_1269), .S(
      n_1268));
   FA_X1 i_635 (.A(p_26[38]), .B(p_27[38]), .CI(p_28[38]), .CO(n_1271), .S(
      n_1270));
   FA_X1 i_636 (.A(p_29[38]), .B(p_30[38]), .CI(n_1223), .CO(n_1273), .S(n_1272));
   FA_X1 i_637 (.A(n_1221), .B(n_1219), .CI(n_1217), .CO(n_1275), .S(n_1274));
   FA_X1 i_638 (.A(n_1215), .B(n_1213), .CI(n_1211), .CO(n_1277), .S(n_1276));
   FA_X1 i_639 (.A(n_1209), .B(n_1931), .CI(n_1229), .CO(n_1279), .S(n_1278));
   FA_X1 i_640 (.A(n_1227), .B(n_1225), .CI(n_1272), .CO(n_1281), .S(n_1280));
   FA_X1 i_641 (.A(n_1270), .B(n_1268), .CI(n_1266), .CO(n_1283), .S(n_1282));
   FA_X1 i_642 (.A(n_1264), .B(n_1262), .CI(n_1260), .CO(n_1285), .S(n_1284));
   FA_X1 i_643 (.A(n_1258), .B(n_1926), .CI(n_1231), .CO(n_1287), .S(n_1286));
   FA_X1 i_644 (.A(n_1278), .B(n_1276), .CI(n_1274), .CO(n_1289), .S(n_1288));
   FA_X1 i_645 (.A(n_1237), .B(n_1235), .CI(n_1233), .CO(n_1291), .S(n_1290));
   FA_X1 i_646 (.A(n_1280), .B(n_1241), .CI(n_1239), .CO(n_1293), .S(n_1292));
   FA_X1 i_647 (.A(n_1286), .B(n_1284), .CI(n_1282), .CO(n_1295), .S(n_1294));
   FA_X1 i_648 (.A(n_1243), .B(n_1290), .CI(n_1288), .CO(n_1297), .S(n_1296));
   FA_X1 i_649 (.A(n_1245), .B(n_1247), .CI(n_1292), .CO(n_1299), .S(n_1298));
   FA_X1 i_650 (.A(n_1249), .B(n_1294), .CI(n_1251), .CO(n_1301), .S(n_1300));
   FA_X1 i_651 (.A(n_1296), .B(n_1298), .CI(n_1253), .CO(n_1303), .S(n_1302));
   FA_X1 i_652 (.A(n_1300), .B(n_1255), .CI(n_1302), .CO(n_1305), .S(n_1304));
   FA_X1 i_653 (.A(p_9[39]), .B(p_10[39]), .CI(p_11[39]), .CO(n_1307), .S(n_1306));
   FA_X1 i_654 (.A(p_12[39]), .B(p_13[39]), .CI(p_14[39]), .CO(n_1309), .S(
      n_1308));
   FA_X1 i_655 (.A(p_15[39]), .B(p_16[39]), .CI(p_17[39]), .CO(n_1311), .S(
      n_1310));
   FA_X1 i_656 (.A(p_18[39]), .B(p_19[39]), .CI(p_20[39]), .CO(n_1313), .S(
      n_1312));
   FA_X1 i_657 (.A(p_21[39]), .B(p_22[39]), .CI(p_23[39]), .CO(n_1315), .S(
      n_1314));
   FA_X1 i_658 (.A(p_24[39]), .B(p_25[39]), .CI(p_26[39]), .CO(n_1317), .S(
      n_1316));
   FA_X1 i_659 (.A(p_27[39]), .B(p_28[39]), .CI(p_29[39]), .CO(n_1319), .S(
      n_1318));
   FA_X1 i_660 (.A(p_30[39]), .B(n_1271), .CI(n_1269), .CO(n_1321), .S(n_1320));
   FA_X1 i_661 (.A(n_1267), .B(n_1265), .CI(n_1263), .CO(n_1323), .S(n_1322));
   FA_X1 i_662 (.A(n_1261), .B(n_1259), .CI(n_1928), .CO(n_1325), .S(n_1324));
   FA_X1 i_663 (.A(n_1277), .B(n_1275), .CI(n_1273), .CO(n_1327), .S(n_1326));
   FA_X1 i_664 (.A(n_1318), .B(n_1316), .CI(n_1314), .CO(n_1329), .S(n_1328));
   FA_X1 i_665 (.A(n_1312), .B(n_1310), .CI(n_1308), .CO(n_1331), .S(n_1330));
   FA_X1 i_666 (.A(n_1306), .B(n_1923), .CI(n_1279), .CO(n_1333), .S(n_1332));
   FA_X1 i_667 (.A(n_1324), .B(n_1322), .CI(n_1320), .CO(n_1335), .S(n_1334));
   FA_X1 i_668 (.A(n_1285), .B(n_1283), .CI(n_1281), .CO(n_1337), .S(n_1336));
   FA_X1 i_669 (.A(n_1287), .B(n_1326), .CI(n_1291), .CO(n_1339), .S(n_1338));
   FA_X1 i_670 (.A(n_1289), .B(n_1332), .CI(n_1330), .CO(n_1341), .S(n_1340));
   FA_X1 i_671 (.A(n_1328), .B(n_1293), .CI(n_1336), .CO(n_1343), .S(n_1342));
   FA_X1 i_672 (.A(n_1334), .B(n_1295), .CI(n_1338), .CO(n_1345), .S(n_1344));
   FA_X1 i_673 (.A(n_1297), .B(n_1340), .CI(n_1342), .CO(n_1347), .S(n_1346));
   FA_X1 i_674 (.A(n_1299), .B(n_1344), .CI(n_1301), .CO(n_1349), .S(n_1348));
   FA_X1 i_675 (.A(n_1303), .B(n_1346), .CI(n_1348), .CO(n_1351), .S(n_1350));
   FA_X1 i_676 (.A(p_10[40]), .B(p_11[40]), .CI(p_12[40]), .CO(n_1353), .S(
      n_1352));
   FA_X1 i_677 (.A(p_13[40]), .B(p_14[40]), .CI(p_15[40]), .CO(n_1355), .S(
      n_1354));
   FA_X1 i_678 (.A(p_16[40]), .B(p_17[40]), .CI(p_18[40]), .CO(n_1357), .S(
      n_1356));
   FA_X1 i_679 (.A(p_19[40]), .B(p_20[40]), .CI(p_21[40]), .CO(n_1359), .S(
      n_1358));
   FA_X1 i_680 (.A(p_22[40]), .B(p_23[40]), .CI(p_24[40]), .CO(n_1361), .S(
      n_1360));
   FA_X1 i_681 (.A(p_25[40]), .B(p_26[40]), .CI(p_27[40]), .CO(n_1363), .S(
      n_1362));
   FA_X1 i_682 (.A(p_28[40]), .B(p_29[40]), .CI(p_30[40]), .CO(n_1365), .S(
      n_1364));
   FA_X1 i_683 (.A(n_1319), .B(n_1317), .CI(n_1315), .CO(n_1367), .S(n_1366));
   FA_X1 i_684 (.A(n_1313), .B(n_1311), .CI(n_1309), .CO(n_1369), .S(n_1368));
   FA_X1 i_685 (.A(n_1307), .B(n_1925), .CI(n_1325), .CO(n_1371), .S(n_1370));
   FA_X1 i_686 (.A(n_1323), .B(n_1321), .CI(n_1364), .CO(n_1373), .S(n_1372));
   FA_X1 i_687 (.A(n_1362), .B(n_1360), .CI(n_1358), .CO(n_1375), .S(n_1374));
   FA_X1 i_688 (.A(n_1356), .B(n_1354), .CI(n_1352), .CO(n_1377), .S(n_1376));
   FA_X1 i_689 (.A(n_1920), .B(n_1327), .CI(n_1370), .CO(n_1379), .S(n_1378));
   FA_X1 i_690 (.A(n_1368), .B(n_1366), .CI(n_1331), .CO(n_1381), .S(n_1380));
   FA_X1 i_691 (.A(n_1329), .B(n_1333), .CI(n_1372), .CO(n_1383), .S(n_1382));
   FA_X1 i_692 (.A(n_1337), .B(n_1335), .CI(n_1376), .CO(n_1385), .S(n_1384));
   FA_X1 i_693 (.A(n_1374), .B(n_1378), .CI(n_1339), .CO(n_1387), .S(n_1386));
   FA_X1 i_694 (.A(n_1380), .B(n_1341), .CI(n_1382), .CO(n_1389), .S(n_1388));
   FA_X1 i_695 (.A(n_1384), .B(n_1343), .CI(n_1386), .CO(n_1391), .S(n_1390));
   FA_X1 i_696 (.A(n_1345), .B(n_1388), .CI(n_1347), .CO(n_1393), .S(n_1392));
   FA_X1 i_697 (.A(n_1390), .B(n_1349), .CI(n_1392), .CO(n_1395), .S(n_1394));
   FA_X1 i_698 (.A(p_11[41]), .B(p_12[41]), .CI(p_13[41]), .CO(n_1397), .S(
      n_1396));
   FA_X1 i_699 (.A(p_14[41]), .B(p_15[41]), .CI(p_16[41]), .CO(n_1399), .S(
      n_1398));
   FA_X1 i_700 (.A(p_17[41]), .B(p_18[41]), .CI(p_19[41]), .CO(n_1401), .S(
      n_1400));
   FA_X1 i_701 (.A(p_20[41]), .B(p_21[41]), .CI(p_22[41]), .CO(n_1403), .S(
      n_1402));
   FA_X1 i_702 (.A(p_23[41]), .B(p_24[41]), .CI(p_25[41]), .CO(n_1405), .S(
      n_1404));
   FA_X1 i_703 (.A(p_26[41]), .B(p_27[41]), .CI(p_28[41]), .CO(n_1407), .S(
      n_1406));
   FA_X1 i_704 (.A(p_29[41]), .B(p_30[41]), .CI(n_1365), .CO(n_1409), .S(n_1408));
   FA_X1 i_705 (.A(n_1363), .B(n_1361), .CI(n_1359), .CO(n_1411), .S(n_1410));
   FA_X1 i_706 (.A(n_1357), .B(n_1355), .CI(n_1353), .CO(n_1413), .S(n_1412));
   FA_X1 i_707 (.A(n_1922), .B(n_1369), .CI(n_1367), .CO(n_1415), .S(n_1414));
   FA_X1 i_708 (.A(n_1408), .B(n_1406), .CI(n_1404), .CO(n_1417), .S(n_1416));
   FA_X1 i_709 (.A(n_1402), .B(n_1400), .CI(n_1398), .CO(n_1419), .S(n_1418));
   FA_X1 i_710 (.A(n_1396), .B(n_1917), .CI(n_1371), .CO(n_1421), .S(n_1420));
   FA_X1 i_711 (.A(n_1412), .B(n_1410), .CI(n_1377), .CO(n_1423), .S(n_1422));
   FA_X1 i_712 (.A(n_1375), .B(n_1373), .CI(n_1414), .CO(n_1425), .S(n_1424));
   FA_X1 i_713 (.A(n_1381), .B(n_1379), .CI(n_1420), .CO(n_1427), .S(n_1426));
   FA_X1 i_714 (.A(n_1418), .B(n_1416), .CI(n_1383), .CO(n_1429), .S(n_1428));
   FA_X1 i_715 (.A(n_1424), .B(n_1422), .CI(n_1385), .CO(n_1431), .S(n_1430));
   FA_X1 i_716 (.A(n_1387), .B(n_1426), .CI(n_1389), .CO(n_1433), .S(n_1432));
   FA_X1 i_717 (.A(n_1428), .B(n_1430), .CI(n_1391), .CO(n_1435), .S(n_1434));
   FA_X1 i_718 (.A(n_1432), .B(n_1393), .CI(n_1434), .CO(n_1437), .S(n_1436));
   FA_X1 i_719 (.A(p_12[42]), .B(p_13[42]), .CI(p_14[42]), .CO(n_1439), .S(
      n_1438));
   FA_X1 i_720 (.A(p_15[42]), .B(p_16[42]), .CI(p_17[42]), .CO(n_1441), .S(
      n_1440));
   FA_X1 i_721 (.A(p_18[42]), .B(p_19[42]), .CI(p_20[42]), .CO(n_1443), .S(
      n_1442));
   FA_X1 i_722 (.A(p_21[42]), .B(p_22[42]), .CI(p_23[42]), .CO(n_1445), .S(
      n_1444));
   FA_X1 i_723 (.A(p_24[42]), .B(p_25[42]), .CI(p_26[42]), .CO(n_1447), .S(
      n_1446));
   FA_X1 i_724 (.A(p_27[42]), .B(p_28[42]), .CI(p_29[42]), .CO(n_1449), .S(
      n_1448));
   FA_X1 i_725 (.A(p_30[42]), .B(n_1407), .CI(n_1405), .CO(n_1451), .S(n_1450));
   FA_X1 i_726 (.A(n_1403), .B(n_1401), .CI(n_1399), .CO(n_1453), .S(n_1452));
   FA_X1 i_727 (.A(n_1397), .B(n_1919), .CI(n_1413), .CO(n_1455), .S(n_1454));
   FA_X1 i_728 (.A(n_1411), .B(n_1409), .CI(n_1448), .CO(n_1457), .S(n_1456));
   FA_X1 i_729 (.A(n_1446), .B(n_1444), .CI(n_1442), .CO(n_1459), .S(n_1458));
   FA_X1 i_730 (.A(n_1440), .B(n_1438), .CI(n_1914), .CO(n_1461), .S(n_1460));
   FA_X1 i_731 (.A(n_1415), .B(n_1454), .CI(n_1452), .CO(n_1463), .S(n_1462));
   FA_X1 i_732 (.A(n_1450), .B(n_1419), .CI(n_1417), .CO(n_1465), .S(n_1464));
   FA_X1 i_733 (.A(n_1421), .B(n_1456), .CI(n_1423), .CO(n_1467), .S(n_1466));
   FA_X1 i_734 (.A(n_1460), .B(n_1458), .CI(n_1425), .CO(n_1469), .S(n_1468));
   FA_X1 i_735 (.A(n_1464), .B(n_1462), .CI(n_1427), .CO(n_1471), .S(n_1470));
   FA_X1 i_736 (.A(n_1429), .B(n_1466), .CI(n_1431), .CO(n_1473), .S(n_1472));
   FA_X1 i_737 (.A(n_1468), .B(n_1433), .CI(n_1470), .CO(n_1475), .S(n_1474));
   FA_X1 i_738 (.A(n_1472), .B(n_1435), .CI(n_1474), .CO(n_1477), .S(n_1476));
   FA_X1 i_739 (.A(p_13[43]), .B(p_14[43]), .CI(p_15[43]), .CO(n_1479), .S(
      n_1478));
   FA_X1 i_740 (.A(p_16[43]), .B(p_17[43]), .CI(p_18[43]), .CO(n_1481), .S(
      n_1480));
   FA_X1 i_741 (.A(p_19[43]), .B(p_20[43]), .CI(p_21[43]), .CO(n_1483), .S(
      n_1482));
   FA_X1 i_742 (.A(p_22[43]), .B(p_23[43]), .CI(p_24[43]), .CO(n_1485), .S(
      n_1484));
   FA_X1 i_743 (.A(p_25[43]), .B(p_26[43]), .CI(p_27[43]), .CO(n_1487), .S(
      n_1486));
   FA_X1 i_744 (.A(p_28[43]), .B(p_29[43]), .CI(p_30[43]), .CO(n_1489), .S(
      n_1488));
   FA_X1 i_745 (.A(n_1449), .B(n_1447), .CI(n_1445), .CO(n_1491), .S(n_1490));
   FA_X1 i_746 (.A(n_1443), .B(n_1441), .CI(n_1439), .CO(n_1493), .S(n_1492));
   FA_X1 i_747 (.A(n_1916), .B(n_1453), .CI(n_1451), .CO(n_1495), .S(n_1494));
   FA_X1 i_748 (.A(n_1488), .B(n_1486), .CI(n_1484), .CO(n_1497), .S(n_1496));
   FA_X1 i_749 (.A(n_1482), .B(n_1480), .CI(n_1478), .CO(n_1499), .S(n_1498));
   FA_X1 i_750 (.A(n_1911), .B(n_1455), .CI(n_1492), .CO(n_1501), .S(n_1500));
   FA_X1 i_751 (.A(n_1490), .B(n_1461), .CI(n_1459), .CO(n_1503), .S(n_1502));
   FA_X1 i_752 (.A(n_1457), .B(n_1494), .CI(n_1465), .CO(n_1505), .S(n_1504));
   FA_X1 i_753 (.A(n_1463), .B(n_1498), .CI(n_1496), .CO(n_1507), .S(n_1506));
   FA_X1 i_754 (.A(n_1500), .B(n_1467), .CI(n_1502), .CO(n_1509), .S(n_1508));
   FA_X1 i_755 (.A(n_1469), .B(n_1504), .CI(n_1471), .CO(n_1511), .S(n_1510));
   FA_X1 i_756 (.A(n_1506), .B(n_1508), .CI(n_1473), .CO(n_1513), .S(n_1512));
   FA_X1 i_757 (.A(n_1510), .B(n_1475), .CI(n_1512), .CO(n_1515), .S(n_1514));
   FA_X1 i_758 (.A(p_14[44]), .B(p_15[44]), .CI(p_16[44]), .CO(n_1517), .S(
      n_1516));
   FA_X1 i_759 (.A(p_17[44]), .B(p_18[44]), .CI(p_19[44]), .CO(n_1519), .S(
      n_1518));
   FA_X1 i_760 (.A(p_20[44]), .B(p_21[44]), .CI(p_22[44]), .CO(n_1521), .S(
      n_1520));
   FA_X1 i_761 (.A(p_23[44]), .B(p_24[44]), .CI(p_25[44]), .CO(n_1523), .S(
      n_1522));
   FA_X1 i_762 (.A(p_26[44]), .B(p_27[44]), .CI(p_28[44]), .CO(n_1525), .S(
      n_1524));
   FA_X1 i_763 (.A(p_29[44]), .B(p_30[44]), .CI(n_1489), .CO(n_1527), .S(n_1526));
   FA_X1 i_764 (.A(n_1487), .B(n_1485), .CI(n_1483), .CO(n_1529), .S(n_1528));
   FA_X1 i_765 (.A(n_1481), .B(n_1479), .CI(n_1913), .CO(n_1531), .S(n_1530));
   FA_X1 i_766 (.A(n_1493), .B(n_1491), .CI(n_1526), .CO(n_1533), .S(n_1532));
   FA_X1 i_767 (.A(n_1524), .B(n_1522), .CI(n_1520), .CO(n_1535), .S(n_1534));
   FA_X1 i_768 (.A(n_1518), .B(n_1516), .CI(n_1908), .CO(n_1537), .S(n_1536));
   FA_X1 i_769 (.A(n_1495), .B(n_1530), .CI(n_1528), .CO(n_1539), .S(n_1538));
   FA_X1 i_770 (.A(n_1499), .B(n_1497), .CI(n_1532), .CO(n_1541), .S(n_1540));
   FA_X1 i_771 (.A(n_1503), .B(n_1501), .CI(n_1536), .CO(n_1543), .S(n_1542));
   FA_X1 i_772 (.A(n_1534), .B(n_1505), .CI(n_1540), .CO(n_1545), .S(n_1544));
   FA_X1 i_773 (.A(n_1538), .B(n_1507), .CI(n_1542), .CO(n_1547), .S(n_1546));
   FA_X1 i_774 (.A(n_1509), .B(n_1544), .CI(n_1511), .CO(n_1549), .S(n_1548));
   FA_X1 i_775 (.A(n_1546), .B(n_1513), .CI(n_1548), .CO(n_1551), .S(n_1550));
   FA_X1 i_776 (.A(p_15[45]), .B(p_16[45]), .CI(p_17[45]), .CO(n_1553), .S(
      n_1552));
   FA_X1 i_777 (.A(p_18[45]), .B(p_19[45]), .CI(p_20[45]), .CO(n_1555), .S(
      n_1554));
   FA_X1 i_778 (.A(p_21[45]), .B(p_22[45]), .CI(p_23[45]), .CO(n_1557), .S(
      n_1556));
   FA_X1 i_779 (.A(p_24[45]), .B(p_25[45]), .CI(p_26[45]), .CO(n_1559), .S(
      n_1558));
   FA_X1 i_780 (.A(p_27[45]), .B(p_28[45]), .CI(p_29[45]), .CO(n_1561), .S(
      n_1560));
   FA_X1 i_781 (.A(p_30[45]), .B(n_1525), .CI(n_1523), .CO(n_1563), .S(n_1562));
   FA_X1 i_782 (.A(n_1521), .B(n_1519), .CI(n_1517), .CO(n_1565), .S(n_1564));
   FA_X1 i_783 (.A(n_1910), .B(n_1531), .CI(n_1529), .CO(n_1567), .S(n_1566));
   FA_X1 i_784 (.A(n_1527), .B(n_1560), .CI(n_1558), .CO(n_1569), .S(n_1568));
   FA_X1 i_785 (.A(n_1556), .B(n_1554), .CI(n_1552), .CO(n_1571), .S(n_1570));
   FA_X1 i_786 (.A(n_1905), .B(n_1564), .CI(n_1562), .CO(n_1573), .S(n_1572));
   FA_X1 i_787 (.A(n_1537), .B(n_1535), .CI(n_1533), .CO(n_1575), .S(n_1574));
   FA_X1 i_788 (.A(n_1566), .B(n_1539), .CI(n_1570), .CO(n_1577), .S(n_1576));
   FA_X1 i_789 (.A(n_1568), .B(n_1541), .CI(n_1574), .CO(n_1579), .S(n_1578));
   FA_X1 i_790 (.A(n_1572), .B(n_1543), .CI(n_1576), .CO(n_1581), .S(n_1580));
   FA_X1 i_791 (.A(n_1545), .B(n_1578), .CI(n_1547), .CO(n_1583), .S(n_1582));
   FA_X1 i_792 (.A(n_1580), .B(n_1549), .CI(n_1582), .CO(n_1585), .S(n_1584));
   FA_X1 i_793 (.A(p_16[46]), .B(p_17[46]), .CI(p_18[46]), .CO(n_1587), .S(
      n_1586));
   FA_X1 i_794 (.A(p_19[46]), .B(p_20[46]), .CI(p_21[46]), .CO(n_1589), .S(
      n_1588));
   FA_X1 i_795 (.A(p_22[46]), .B(p_23[46]), .CI(p_24[46]), .CO(n_1591), .S(
      n_1590));
   FA_X1 i_796 (.A(p_25[46]), .B(p_26[46]), .CI(p_27[46]), .CO(n_1593), .S(
      n_1592));
   FA_X1 i_797 (.A(p_28[46]), .B(p_29[46]), .CI(p_30[46]), .CO(n_1595), .S(
      n_1594));
   FA_X1 i_798 (.A(n_1561), .B(n_1559), .CI(n_1557), .CO(n_1597), .S(n_1596));
   FA_X1 i_799 (.A(n_1555), .B(n_1553), .CI(n_1907), .CO(n_1599), .S(n_1598));
   FA_X1 i_800 (.A(n_1565), .B(n_1563), .CI(n_1594), .CO(n_1601), .S(n_1600));
   FA_X1 i_801 (.A(n_1592), .B(n_1590), .CI(n_1588), .CO(n_1603), .S(n_1602));
   FA_X1 i_802 (.A(n_1586), .B(n_1902), .CI(n_1567), .CO(n_1605), .S(n_1604));
   FA_X1 i_803 (.A(n_1598), .B(n_1596), .CI(n_1571), .CO(n_1607), .S(n_1606));
   FA_X1 i_804 (.A(n_1569), .B(n_1600), .CI(n_1575), .CO(n_1609), .S(n_1608));
   FA_X1 i_805 (.A(n_1573), .B(n_1604), .CI(n_1602), .CO(n_1611), .S(n_1610));
   FA_X1 i_806 (.A(n_1606), .B(n_1577), .CI(n_1608), .CO(n_1613), .S(n_1612));
   FA_X1 i_807 (.A(n_1579), .B(n_1610), .CI(n_1581), .CO(n_1615), .S(n_1614));
   FA_X1 i_808 (.A(n_1612), .B(n_1583), .CI(n_1614), .CO(n_1617), .S(n_1616));
   FA_X1 i_809 (.A(p_17[47]), .B(p_18[47]), .CI(p_19[47]), .CO(n_1619), .S(
      n_1618));
   FA_X1 i_810 (.A(p_20[47]), .B(p_21[47]), .CI(p_22[47]), .CO(n_1621), .S(
      n_1620));
   FA_X1 i_811 (.A(p_23[47]), .B(p_24[47]), .CI(p_25[47]), .CO(n_1623), .S(
      n_1622));
   FA_X1 i_812 (.A(p_26[47]), .B(p_27[47]), .CI(p_28[47]), .CO(n_1625), .S(
      n_1624));
   FA_X1 i_813 (.A(p_29[47]), .B(p_30[47]), .CI(n_1595), .CO(n_1627), .S(n_1626));
   FA_X1 i_814 (.A(n_1593), .B(n_1591), .CI(n_1589), .CO(n_1629), .S(n_1628));
   FA_X1 i_815 (.A(n_1587), .B(n_1904), .CI(n_1599), .CO(n_1631), .S(n_1630));
   FA_X1 i_816 (.A(n_1597), .B(n_1626), .CI(n_1624), .CO(n_1633), .S(n_1632));
   FA_X1 i_817 (.A(n_1622), .B(n_1620), .CI(n_1618), .CO(n_1635), .S(n_1634));
   FA_X1 i_818 (.A(n_1899), .B(n_1630), .CI(n_1628), .CO(n_1637), .S(n_1636));
   FA_X1 i_819 (.A(n_1603), .B(n_1601), .CI(n_1605), .CO(n_1639), .S(n_1638));
   FA_X1 i_820 (.A(n_1607), .B(n_1634), .CI(n_1632), .CO(n_1641), .S(n_1640));
   FA_X1 i_821 (.A(n_1609), .B(n_1638), .CI(n_1636), .CO(n_1643), .S(n_1642));
   FA_X1 i_822 (.A(n_1611), .B(n_1640), .CI(n_1613), .CO(n_1645), .S(n_1644));
   FA_X1 i_823 (.A(n_1642), .B(n_1615), .CI(n_1644), .CO(n_1647), .S(n_1646));
   FA_X1 i_824 (.A(p_18[48]), .B(p_19[48]), .CI(p_20[48]), .CO(n_1649), .S(
      n_1648));
   FA_X1 i_825 (.A(p_21[48]), .B(p_22[48]), .CI(p_23[48]), .CO(n_1651), .S(
      n_1650));
   FA_X1 i_826 (.A(p_24[48]), .B(p_25[48]), .CI(p_26[48]), .CO(n_1653), .S(
      n_1652));
   FA_X1 i_827 (.A(p_27[48]), .B(p_28[48]), .CI(p_29[48]), .CO(n_1655), .S(
      n_1654));
   FA_X1 i_828 (.A(p_30[48]), .B(n_1625), .CI(n_1623), .CO(n_1657), .S(n_1656));
   FA_X1 i_829 (.A(n_1621), .B(n_1619), .CI(n_1901), .CO(n_1659), .S(n_1658));
   FA_X1 i_830 (.A(n_1629), .B(n_1627), .CI(n_1654), .CO(n_1661), .S(n_1660));
   FA_X1 i_831 (.A(n_1652), .B(n_1650), .CI(n_1648), .CO(n_1663), .S(n_1662));
   FA_X1 i_832 (.A(n_1896), .B(n_1631), .CI(n_1658), .CO(n_1665), .S(n_1664));
   FA_X1 i_833 (.A(n_1656), .B(n_1635), .CI(n_1633), .CO(n_1667), .S(n_1666));
   FA_X1 i_834 (.A(n_1660), .B(n_1637), .CI(n_1639), .CO(n_1669), .S(n_1668));
   FA_X1 i_835 (.A(n_1662), .B(n_1664), .CI(n_1666), .CO(n_1671), .S(n_1670));
   FA_X1 i_836 (.A(n_1641), .B(n_1668), .CI(n_1643), .CO(n_1673), .S(n_1672));
   FA_X1 i_837 (.A(n_1670), .B(n_1645), .CI(n_1672), .CO(n_1675), .S(n_1674));
   FA_X1 i_838 (.A(p_19[49]), .B(p_20[49]), .CI(p_21[49]), .CO(n_1677), .S(
      n_1676));
   FA_X1 i_839 (.A(p_22[49]), .B(p_23[49]), .CI(p_24[49]), .CO(n_1679), .S(
      n_1678));
   FA_X1 i_840 (.A(p_25[49]), .B(p_26[49]), .CI(p_27[49]), .CO(n_1681), .S(
      n_1680));
   FA_X1 i_841 (.A(p_28[49]), .B(p_29[49]), .CI(p_30[49]), .CO(n_1683), .S(
      n_1682));
   FA_X1 i_842 (.A(n_1655), .B(n_1653), .CI(n_1651), .CO(n_1685), .S(n_1684));
   FA_X1 i_843 (.A(n_1649), .B(n_1898), .CI(n_1659), .CO(n_1687), .S(n_1686));
   FA_X1 i_844 (.A(n_1657), .B(n_1682), .CI(n_1680), .CO(n_1689), .S(n_1688));
   FA_X1 i_845 (.A(n_1678), .B(n_1676), .CI(n_1893), .CO(n_1691), .S(n_1690));
   FA_X1 i_846 (.A(n_1686), .B(n_1684), .CI(n_1663), .CO(n_1693), .S(n_1692));
   FA_X1 i_847 (.A(n_1661), .B(n_1667), .CI(n_1665), .CO(n_1695), .S(n_1694));
   FA_X1 i_848 (.A(n_1690), .B(n_1688), .CI(n_1669), .CO(n_1697), .S(n_1696));
   FA_X1 i_849 (.A(n_1692), .B(n_1694), .CI(n_1671), .CO(n_1699), .S(n_1698));
   FA_X1 i_850 (.A(n_1696), .B(n_1673), .CI(n_1698), .CO(n_1701), .S(n_1700));
   FA_X1 i_851 (.A(p_20[50]), .B(p_21[50]), .CI(p_22[50]), .CO(n_1703), .S(
      n_1702));
   FA_X1 i_852 (.A(p_23[50]), .B(p_24[50]), .CI(p_25[50]), .CO(n_1705), .S(
      n_1704));
   FA_X1 i_853 (.A(p_26[50]), .B(p_27[50]), .CI(p_28[50]), .CO(n_1707), .S(
      n_1706));
   FA_X1 i_854 (.A(p_29[50]), .B(p_30[50]), .CI(n_1683), .CO(n_1709), .S(n_1708));
   FA_X1 i_855 (.A(n_1681), .B(n_1679), .CI(n_1677), .CO(n_1711), .S(n_1710));
   FA_X1 i_856 (.A(n_1895), .B(n_1685), .CI(n_1708), .CO(n_1713), .S(n_1712));
   FA_X1 i_857 (.A(n_1706), .B(n_1704), .CI(n_1702), .CO(n_1715), .S(n_1714));
   FA_X1 i_858 (.A(n_1890), .B(n_1687), .CI(n_1710), .CO(n_1717), .S(n_1716));
   FA_X1 i_859 (.A(n_1691), .B(n_1689), .CI(n_1712), .CO(n_1719), .S(n_1718));
   FA_X1 i_860 (.A(n_1693), .B(n_1714), .CI(n_1716), .CO(n_1721), .S(n_1720));
   FA_X1 i_861 (.A(n_1695), .B(n_1718), .CI(n_1697), .CO(n_1723), .S(n_1722));
   FA_X1 i_862 (.A(n_1720), .B(n_1699), .CI(n_1722), .CO(n_1725), .S(n_1724));
   FA_X1 i_863 (.A(p_21[51]), .B(p_22[51]), .CI(p_23[51]), .CO(n_1727), .S(
      n_1726));
   FA_X1 i_864 (.A(p_24[51]), .B(p_25[51]), .CI(p_26[51]), .CO(n_1729), .S(
      n_1728));
   FA_X1 i_865 (.A(p_27[51]), .B(p_28[51]), .CI(p_29[51]), .CO(n_1731), .S(
      n_1730));
   FA_X1 i_866 (.A(p_30[51]), .B(n_1707), .CI(n_1705), .CO(n_1733), .S(n_1732));
   FA_X1 i_867 (.A(n_1703), .B(n_1892), .CI(n_1711), .CO(n_1735), .S(n_1734));
   FA_X1 i_868 (.A(n_1709), .B(n_1730), .CI(n_1728), .CO(n_1737), .S(n_1736));
   FA_X1 i_869 (.A(n_1726), .B(n_1887), .CI(n_1734), .CO(n_1739), .S(n_1738));
   FA_X1 i_870 (.A(n_1732), .B(n_1715), .CI(n_1713), .CO(n_1741), .S(n_1740));
   FA_X1 i_871 (.A(n_1717), .B(n_1738), .CI(n_1736), .CO(n_1743), .S(n_1742));
   FA_X1 i_872 (.A(n_1719), .B(n_1740), .CI(n_1721), .CO(n_1745), .S(n_1744));
   FA_X1 i_873 (.A(n_1723), .B(n_1742), .CI(n_1744), .CO(n_1747), .S(n_1746));
   FA_X1 i_874 (.A(p_22[52]), .B(p_23[52]), .CI(p_24[52]), .CO(n_1749), .S(
      n_1748));
   FA_X1 i_875 (.A(p_25[52]), .B(p_26[52]), .CI(p_27[52]), .CO(n_1751), .S(
      n_1750));
   FA_X1 i_876 (.A(p_28[52]), .B(p_29[52]), .CI(p_30[52]), .CO(n_1753), .S(
      n_1752));
   FA_X1 i_877 (.A(n_1731), .B(n_1729), .CI(n_1727), .CO(n_1755), .S(n_1754));
   FA_X1 i_878 (.A(n_1889), .B(n_1733), .CI(n_1752), .CO(n_1757), .S(n_1756));
   FA_X1 i_879 (.A(n_1750), .B(n_1748), .CI(n_1884), .CO(n_1759), .S(n_1758));
   FA_X1 i_880 (.A(n_1735), .B(n_1754), .CI(n_1737), .CO(n_1761), .S(n_1760));
   FA_X1 i_881 (.A(n_1756), .B(n_1741), .CI(n_1739), .CO(n_1763), .S(n_1762));
   FA_X1 i_882 (.A(n_1758), .B(n_1760), .CI(n_1743), .CO(n_1765), .S(n_1764));
   FA_X1 i_883 (.A(n_1762), .B(n_1745), .CI(n_1764), .CO(n_1767), .S(n_1766));
   FA_X1 i_884 (.A(p_23[53]), .B(p_24[53]), .CI(p_25[53]), .CO(n_1769), .S(
      n_1768));
   FA_X1 i_885 (.A(p_26[53]), .B(p_27[53]), .CI(p_28[53]), .CO(n_1771), .S(
      n_1770));
   FA_X1 i_886 (.A(p_29[53]), .B(p_30[53]), .CI(n_1753), .CO(n_1773), .S(n_1772));
   FA_X1 i_887 (.A(n_1751), .B(n_1749), .CI(n_1886), .CO(n_1775), .S(n_1774));
   FA_X1 i_888 (.A(n_1755), .B(n_1772), .CI(n_1770), .CO(n_1777), .S(n_1776));
   FA_X1 i_889 (.A(n_1768), .B(n_1881), .CI(n_1774), .CO(n_1779), .S(n_1778));
   FA_X1 i_890 (.A(n_1759), .B(n_1757), .CI(n_1761), .CO(n_1781), .S(n_1780));
   FA_X1 i_891 (.A(n_1778), .B(n_1776), .CI(n_1763), .CO(n_1783), .S(n_1782));
   FA_X1 i_892 (.A(n_1780), .B(n_1765), .CI(n_1782), .CO(n_1785), .S(n_1784));
   FA_X1 i_893 (.A(p_24[54]), .B(p_25[54]), .CI(p_26[54]), .CO(n_1787), .S(
      n_1786));
   FA_X1 i_894 (.A(p_27[54]), .B(p_28[54]), .CI(p_29[54]), .CO(n_1789), .S(
      n_1788));
   FA_X1 i_895 (.A(p_30[54]), .B(n_1771), .CI(n_1769), .CO(n_1791), .S(n_1790));
   FA_X1 i_896 (.A(n_1883), .B(n_1775), .CI(n_1773), .CO(n_1793), .S(n_1792));
   FA_X1 i_897 (.A(n_1788), .B(n_1786), .CI(n_1878), .CO(n_1795), .S(n_1794));
   FA_X1 i_898 (.A(n_1790), .B(n_1777), .CI(n_1792), .CO(n_1797), .S(n_1796));
   FA_X1 i_899 (.A(n_1779), .B(n_1794), .CI(n_1781), .CO(n_1799), .S(n_1798));
   FA_X1 i_900 (.A(n_1796), .B(n_1783), .CI(n_1798), .CO(n_1801), .S(n_1800));
   FA_X1 i_901 (.A(p_25[55]), .B(p_26[55]), .CI(p_27[55]), .CO(n_1803), .S(
      n_1802));
   FA_X1 i_902 (.A(p_28[55]), .B(p_29[55]), .CI(p_30[55]), .CO(n_1805), .S(
      n_1804));
   FA_X1 i_903 (.A(n_1789), .B(n_1787), .CI(n_1880), .CO(n_1807), .S(n_1806));
   FA_X1 i_904 (.A(n_1791), .B(n_1804), .CI(n_1802), .CO(n_1809), .S(n_1808));
   FA_X1 i_905 (.A(n_1875), .B(n_1793), .CI(n_1806), .CO(n_1811), .S(n_1810));
   FA_X1 i_906 (.A(n_1795), .B(n_1808), .CI(n_1810), .CO(n_1813), .S(n_1812));
   FA_X1 i_907 (.A(n_1797), .B(n_1799), .CI(n_1812), .CO(n_1815), .S(n_1814));
   FA_X1 i_908 (.A(p_26[56]), .B(p_27[56]), .CI(p_28[56]), .CO(n_1817), .S(
      n_1816));
   FA_X1 i_909 (.A(p_29[56]), .B(p_30[56]), .CI(n_1805), .CO(n_1819), .S(n_1818));
   FA_X1 i_910 (.A(n_1803), .B(n_1877), .CI(n_1807), .CO(n_1821), .S(n_1820));
   FA_X1 i_911 (.A(n_1818), .B(n_1816), .CI(n_1872), .CO(n_1823), .S(n_1822));
   FA_X1 i_912 (.A(n_1820), .B(n_1809), .CI(n_1811), .CO(n_1825), .S(n_1824));
   FA_X1 i_913 (.A(n_1822), .B(n_1824), .CI(n_1813), .CO(n_1827), .S(n_1826));
   FA_X1 i_914 (.A(p_27[57]), .B(p_28[57]), .CI(p_29[57]), .CO(n_1829), .S(
      n_1828));
   FA_X1 i_915 (.A(p_30[57]), .B(n_1817), .CI(n_1874), .CO(n_1831), .S(n_1830));
   FA_X1 i_916 (.A(n_1819), .B(n_1828), .CI(n_1869), .CO(n_1833), .S(n_1832));
   FA_X1 i_917 (.A(n_1821), .B(n_1830), .CI(n_1823), .CO(n_1835), .S(n_1834));
   FA_X1 i_918 (.A(n_1832), .B(n_1825), .CI(n_1834), .CO(n_1837), .S(n_1836));
   FA_X1 i_919 (.A(p_28[58]), .B(p_29[58]), .CI(p_30[58]), .CO(n_1839), .S(
      n_1838));
   FA_X1 i_920 (.A(n_1829), .B(n_1871), .CI(n_1831), .CO(n_1841), .S(n_1840));
   FA_X1 i_921 (.A(n_1838), .B(n_1866), .CI(n_1840), .CO(n_1843), .S(n_1842));
   FA_X1 i_922 (.A(n_1833), .B(n_1835), .CI(n_1842), .CO(n_1845), .S(n_1844));
   FA_X1 i_923 (.A(p_29[59]), .B(p_30[59]), .CI(n_1839), .CO(n_1847), .S(n_1846));
   FA_X1 i_924 (.A(n_1868), .B(n_1846), .CI(n_1863), .CO(n_1849), .S(n_1848));
   FA_X1 i_925 (.A(n_1841), .B(n_1843), .CI(n_1848), .CO(n_1851), .S(n_1850));
   FA_X1 i_926 (.A(p_30[60]), .B(n_1865), .CI(n_1847), .CO(n_1853), .S(n_1852));
   FA_X1 i_927 (.A(n_1860), .B(n_1852), .CI(n_1849), .CO(n_1855), .S(n_1854));
   FA_X1 i_928 (.A(n_1862), .B(n_1858), .CI(n_1853), .CO(n_1857), .S(n_1856));
   XNOR2_X1 i_929 (.A(p_29[61]), .B(n_1859), .ZN(n_1858));
   OAI21_X1 i_930 (.A(n_2322), .B1(n_2335), .B2(p_30[61]), .ZN(n_1859));
   XOR2_X1 i_931 (.A(n_2332), .B(n_1861), .Z(n_1860));
   XOR2_X1 i_932 (.A(p_27[60]), .B(p_28[60]), .Z(n_1861));
   OAI222_X1 i_933 (.A1(p_27[60]), .A2(n_2332), .B1(p_27[60]), .B2(n_2334), 
      .C1(n_2334), .C2(n_2332), .ZN(n_1862));
   XOR2_X1 i_934 (.A(n_2333), .B(n_1864), .Z(n_1863));
   XOR2_X1 i_935 (.A(p_26[62]), .B(p_27[59]), .Z(n_1864));
   OAI222_X1 i_936 (.A1(p_26[62]), .A2(n_2333), .B1(p_26[62]), .B2(n_2337), 
      .C1(n_2337), .C2(n_2333), .ZN(n_1865));
   XOR2_X1 i_937 (.A(n_2336), .B(n_1867), .Z(n_1866));
   XOR2_X1 i_938 (.A(p_25[62]), .B(p_26[58]), .Z(n_1867));
   OAI222_X1 i_939 (.A1(p_25[62]), .A2(n_2336), .B1(p_25[62]), .B2(n_2339), 
      .C1(n_2339), .C2(n_2336), .ZN(n_1868));
   XOR2_X1 i_940 (.A(n_2338), .B(n_1870), .Z(n_1869));
   XOR2_X1 i_941 (.A(p_24[62]), .B(p_25[57]), .Z(n_1870));
   OAI222_X1 i_942 (.A1(p_24[62]), .A2(n_2338), .B1(p_24[62]), .B2(n_2341), 
      .C1(n_2341), .C2(n_2338), .ZN(n_1871));
   XOR2_X1 i_943 (.A(n_2340), .B(n_1873), .Z(n_1872));
   XOR2_X1 i_944 (.A(p_23[62]), .B(p_24[56]), .Z(n_1873));
   OAI222_X1 i_945 (.A1(p_23[62]), .A2(n_2340), .B1(p_23[62]), .B2(n_2343), 
      .C1(n_2343), .C2(n_2340), .ZN(n_1874));
   XOR2_X1 i_946 (.A(n_2342), .B(n_1876), .Z(n_1875));
   XOR2_X1 i_947 (.A(p_22[62]), .B(p_23[55]), .Z(n_1876));
   OAI222_X1 i_948 (.A1(p_22[62]), .A2(n_2342), .B1(p_22[62]), .B2(n_2345), 
      .C1(n_2345), .C2(n_2342), .ZN(n_1877));
   XOR2_X1 i_949 (.A(n_2344), .B(n_1879), .Z(n_1878));
   XOR2_X1 i_950 (.A(p_21[62]), .B(p_22[54]), .Z(n_1879));
   OAI222_X1 i_951 (.A1(p_21[62]), .A2(n_2344), .B1(p_21[62]), .B2(n_2347), 
      .C1(n_2347), .C2(n_2344), .ZN(n_1880));
   XOR2_X1 i_952 (.A(n_2346), .B(n_1882), .Z(n_1881));
   XOR2_X1 i_953 (.A(p_20[62]), .B(p_21[53]), .Z(n_1882));
   OAI222_X1 i_954 (.A1(p_20[62]), .A2(n_2346), .B1(p_20[62]), .B2(n_2349), 
      .C1(n_2349), .C2(n_2346), .ZN(n_1883));
   XOR2_X1 i_955 (.A(n_2348), .B(n_1885), .Z(n_1884));
   XOR2_X1 i_956 (.A(p_19[62]), .B(p_20[52]), .Z(n_1885));
   OAI222_X1 i_957 (.A1(p_19[62]), .A2(n_2348), .B1(p_19[62]), .B2(n_2351), 
      .C1(n_2351), .C2(n_2348), .ZN(n_1886));
   XOR2_X1 i_958 (.A(n_2350), .B(n_1888), .Z(n_1887));
   XOR2_X1 i_959 (.A(p_18[62]), .B(p_19[51]), .Z(n_1888));
   OAI222_X1 i_960 (.A1(p_18[62]), .A2(n_2350), .B1(p_18[62]), .B2(n_2353), 
      .C1(n_2353), .C2(n_2350), .ZN(n_1889));
   XOR2_X1 i_961 (.A(n_2352), .B(n_1891), .Z(n_1890));
   XOR2_X1 i_962 (.A(p_17[62]), .B(p_18[50]), .Z(n_1891));
   OAI222_X1 i_963 (.A1(p_17[62]), .A2(n_2352), .B1(p_17[62]), .B2(n_2355), 
      .C1(n_2355), .C2(n_2352), .ZN(n_1892));
   XOR2_X1 i_964 (.A(n_2354), .B(n_1894), .Z(n_1893));
   XOR2_X1 i_965 (.A(p_16[62]), .B(p_17[49]), .Z(n_1894));
   OAI222_X1 i_966 (.A1(p_16[62]), .A2(n_2354), .B1(p_16[62]), .B2(n_2357), 
      .C1(n_2357), .C2(n_2354), .ZN(n_1895));
   XOR2_X1 i_967 (.A(n_2356), .B(n_1897), .Z(n_1896));
   XOR2_X1 i_968 (.A(p_15[62]), .B(p_16[48]), .Z(n_1897));
   OAI222_X1 i_969 (.A1(p_15[62]), .A2(n_2356), .B1(p_15[62]), .B2(n_2359), 
      .C1(n_2359), .C2(n_2356), .ZN(n_1898));
   XOR2_X1 i_970 (.A(n_2358), .B(n_1900), .Z(n_1899));
   XOR2_X1 i_971 (.A(p_14[62]), .B(p_15[47]), .Z(n_1900));
   OAI222_X1 i_972 (.A1(p_14[62]), .A2(n_2358), .B1(p_14[62]), .B2(n_2361), 
      .C1(n_2361), .C2(n_2358), .ZN(n_1901));
   XOR2_X1 i_973 (.A(n_2360), .B(n_1903), .Z(n_1902));
   XOR2_X1 i_974 (.A(p_13[62]), .B(p_14[46]), .Z(n_1903));
   OAI222_X1 i_975 (.A1(p_13[62]), .A2(n_2360), .B1(p_13[62]), .B2(n_2363), 
      .C1(n_2363), .C2(n_2360), .ZN(n_1904));
   XOR2_X1 i_976 (.A(n_2362), .B(n_1906), .Z(n_1905));
   XOR2_X1 i_977 (.A(p_12[62]), .B(p_13[45]), .Z(n_1906));
   OAI222_X1 i_978 (.A1(p_12[62]), .A2(n_2362), .B1(p_12[62]), .B2(n_2365), 
      .C1(n_2365), .C2(n_2362), .ZN(n_1907));
   XOR2_X1 i_979 (.A(n_2364), .B(n_1909), .Z(n_1908));
   XOR2_X1 i_980 (.A(p_11[62]), .B(p_12[44]), .Z(n_1909));
   OAI222_X1 i_981 (.A1(p_11[62]), .A2(n_2364), .B1(p_11[62]), .B2(n_2367), 
      .C1(n_2367), .C2(n_2364), .ZN(n_1910));
   XOR2_X1 i_982 (.A(n_2366), .B(n_1912), .Z(n_1911));
   XOR2_X1 i_983 (.A(p_10[62]), .B(p_11[43]), .Z(n_1912));
   OAI222_X1 i_984 (.A1(p_10[62]), .A2(n_2366), .B1(p_10[62]), .B2(n_2369), 
      .C1(n_2369), .C2(n_2366), .ZN(n_1913));
   XOR2_X1 i_985 (.A(n_2368), .B(n_1915), .Z(n_1914));
   XOR2_X1 i_986 (.A(p_9[62]), .B(p_10[42]), .Z(n_1915));
   OAI222_X1 i_987 (.A1(p_9[62]), .A2(n_2368), .B1(p_9[62]), .B2(n_2371), 
      .C1(n_2371), .C2(n_2368), .ZN(n_1916));
   XOR2_X1 i_988 (.A(n_2370), .B(n_1918), .Z(n_1917));
   XOR2_X1 i_989 (.A(p_8[59]), .B(p_9[41]), .Z(n_1918));
   OAI222_X1 i_990 (.A1(p_8[59]), .A2(n_2370), .B1(p_8[59]), .B2(n_2373), 
      .C1(n_2373), .C2(n_2370), .ZN(n_1919));
   XOR2_X1 i_991 (.A(n_2372), .B(n_1921), .Z(n_1920));
   XOR2_X1 i_992 (.A(p_7[59]), .B(p_8[40]), .Z(n_1921));
   OAI222_X1 i_993 (.A1(p_7[59]), .A2(n_2372), .B1(p_7[59]), .B2(n_2375), 
      .C1(n_2375), .C2(n_2372), .ZN(n_1922));
   XOR2_X1 i_997 (.A(n_2376), .B(n_1927), .Z(n_1926));
   XOR2_X1 i_998 (.A(p_5[59]), .B(p_6[38]), .Z(n_1927));
   XOR2_X1 i_1003 (.A(n_2380), .B(n_1933), .Z(n_1932));
   XOR2_X1 i_1004 (.A(p_3[59]), .B(p_4[36]), .Z(n_1933));
   XOR2_X1 i_1006 (.A(n_2382), .B(n_1936), .Z(n_1935));
   XOR2_X1 i_1007 (.A(p_2[59]), .B(p_3[35]), .Z(n_1936));
   OAI222_X1 i_1008 (.A1(p_2[59]), .A2(n_2382), .B1(p_2[59]), .B2(n_2385), 
      .C1(n_2385), .C2(n_2382), .ZN(n_1937));
   OAI222_X1 i_1014 (.A1(p_0[59]), .A2(n_2386), .B1(p_0[59]), .B2(n_2389), 
      .C1(n_2389), .C2(n_2386), .ZN(n_1943));
   AOI22_X1 i_1015 (.A1(out[61]), .A2(n_1945), .B1(n_1947), .B2(n_1946), 
      .ZN(n_1944));
   OAI21_X1 i_1016 (.A(n_1947), .B1(p_29[32]), .B2(p_30[32]), .ZN(n_1945));
   OAI21_X1 i_1020 (.A(n_1950), .B1(n_2390), .B2(n_2388), .ZN(n_1949));
   NAND2_X1 i_1021 (.A1(n_2390), .A2(n_2388), .ZN(n_1950));
   INV_X1 i_1022 (.A(n_1951), .ZN(out31[1]));
   OAI21_X1 i_1023 (.A(n_2310), .B1(p_0[1]), .B2(out[1]), .ZN(n_1951));
   XOR2_X1 i_1024 (.A(n_2310), .B(n_1952), .Z(out31[2]));
   OAI21_X1 i_1025 (.A(n_2309), .B1(out[2]), .B2(n_0), .ZN(n_1952));
   XNOR2_X1 i_1026 (.A(n_2308), .B(n_1953), .ZN(out31[3]));
   OAI21_X1 i_1027 (.A(n_2313), .B1(n_2), .B2(n_4), .ZN(n_1953));
   XOR2_X1 i_1028 (.A(n_2307), .B(n_1954), .Z(out31[4]));
   OAI21_X1 i_1029 (.A(n_2314), .B1(n_2330), .B2(n_2329), .ZN(n_1954));
   XOR2_X1 i_1030 (.A(n_2305), .B(n_1961), .Z(out31[5]));
   XOR2_X1 i_1031 (.A(n_1960), .B(n_1957), .Z(out31[6]));
   XOR2_X1 i_1032 (.A(n_1958), .B(n_1955), .Z(out31[7]));
   NOR2_X1 i_1033 (.A1(n_2302), .A2(n_2293), .ZN(n_1955));
   XNOR2_X1 i_1034 (.A(n_1962), .B(n_1956), .ZN(out31[8]));
   OAI22_X1 i_1035 (.A1(n_38), .A2(n_40), .B1(n_2293), .B2(n_1958), .ZN(n_1956));
   AOI21_X1 i_1036 (.A(n_2303), .B1(n_26), .B2(n_28), .ZN(n_1957));
   AOI21_X1 i_1037 (.A(n_2303), .B1(n_2297), .B2(n_1959), .ZN(n_1958));
   INV_X1 i_1038 (.A(n_1960), .ZN(n_1959));
   AOI21_X1 i_1039 (.A(n_2300), .B1(n_2305), .B2(n_2298), .ZN(n_1960));
   OAI21_X1 i_1040 (.A(n_2298), .B1(n_16), .B2(n_18), .ZN(n_1961));
   NOR2_X1 i_1041 (.A1(n_2304), .A2(n_2295), .ZN(n_1962));
   XNOR2_X1 i_1042 (.A(n_2291), .B(n_1969), .ZN(out31[9]));
   XOR2_X1 i_1043 (.A(n_1968), .B(n_1965), .Z(out31[10]));
   XOR2_X1 i_1044 (.A(n_1966), .B(n_1963), .Z(out31[11]));
   NOR2_X1 i_1045 (.A1(n_2288), .A2(n_2279), .ZN(n_1963));
   XNOR2_X1 i_1046 (.A(n_1970), .B(n_1964), .ZN(out31[12]));
   OAI22_X1 i_1047 (.A1(n_106), .A2(n_108), .B1(n_2279), .B2(n_1966), .ZN(n_1964));
   AOI21_X1 i_1048 (.A(n_2289), .B1(n_86), .B2(n_88), .ZN(n_1965));
   AOI21_X1 i_1049 (.A(n_2289), .B1(n_2283), .B2(n_1967), .ZN(n_1966));
   INV_X1 i_1050 (.A(n_1968), .ZN(n_1967));
   AOI21_X1 i_1051 (.A(n_2286), .B1(n_2291), .B2(n_2284), .ZN(n_1968));
   AOI21_X1 i_1052 (.A(n_2286), .B1(n_68), .B2(n_70), .ZN(n_1969));
   NOR2_X1 i_1053 (.A1(n_2290), .A2(n_2281), .ZN(n_1970));
   XOR2_X1 i_1054 (.A(n_2277), .B(n_1977), .Z(out31[13]));
   XOR2_X1 i_1055 (.A(n_1976), .B(n_1973), .Z(out31[14]));
   XOR2_X1 i_1056 (.A(n_1974), .B(n_1971), .Z(out31[15]));
   NOR2_X1 i_1057 (.A1(n_2274), .A2(n_2265), .ZN(n_1971));
   XNOR2_X1 i_1058 (.A(n_1978), .B(n_1972), .ZN(out31[16]));
   OAI22_X1 i_1059 (.A1(n_206), .A2(n_208), .B1(n_2265), .B2(n_1974), .ZN(n_1972));
   AOI21_X1 i_1060 (.A(n_2275), .B1(n_178), .B2(n_180), .ZN(n_1973));
   AOI21_X1 i_1061 (.A(n_2275), .B1(n_2269), .B2(n_1975), .ZN(n_1974));
   INV_X1 i_1062 (.A(n_1976), .ZN(n_1975));
   AOI21_X1 i_1063 (.A(n_2272), .B1(n_2277), .B2(n_2270), .ZN(n_1976));
   OAI21_X1 i_1064 (.A(n_2270), .B1(n_152), .B2(n_154), .ZN(n_1977));
   NOR2_X1 i_1065 (.A1(n_2276), .A2(n_2267), .ZN(n_1978));
   XOR2_X1 i_1066 (.A(n_2263), .B(n_1985), .Z(out31[17]));
   XOR2_X1 i_1067 (.A(n_1984), .B(n_1981), .Z(out31[18]));
   XOR2_X1 i_1068 (.A(n_1982), .B(n_1979), .Z(out31[19]));
   NOR2_X1 i_1069 (.A1(n_2229), .A2(n_2219), .ZN(n_1979));
   XNOR2_X1 i_1070 (.A(n_1986), .B(n_1980), .ZN(out31[20]));
   OAI21_X1 i_1071 (.A(n_2228), .B1(n_2219), .B2(n_1982), .ZN(n_1980));
   NOR2_X1 i_1072 (.A1(n_2231), .A2(n_2221), .ZN(n_1981));
   INV_X1 i_1073 (.A(n_1983), .ZN(n_1982));
   OAI21_X1 i_1074 (.A(n_2230), .B1(n_2221), .B2(n_1984), .ZN(n_1983));
   AOI21_X1 i_1075 (.A(n_2226), .B1(n_2263), .B2(n_2223), .ZN(n_1984));
   OAI21_X1 i_1076 (.A(n_2223), .B1(n_268), .B2(n_270), .ZN(n_1985));
   AOI21_X1 i_1077 (.A(n_2233), .B1(n_376), .B2(n_378), .ZN(n_1986));
   XOR2_X1 i_1078 (.A(n_2014), .B(n_1993), .Z(out31[21]));
   XOR2_X1 i_1079 (.A(n_1992), .B(n_1989), .Z(out31[22]));
   XOR2_X1 i_1080 (.A(n_1990), .B(n_1987), .Z(out31[23]));
   NOR2_X1 i_1081 (.A1(n_2257), .A2(n_2201), .ZN(n_1987));
   XNOR2_X1 i_1082 (.A(n_1994), .B(n_1988), .ZN(out31[24]));
   OAI21_X1 i_1083 (.A(n_2256), .B1(n_2201), .B2(n_1990), .ZN(n_1988));
   NOR2_X1 i_1084 (.A1(n_2259), .A2(n_2203), .ZN(n_1989));
   INV_X1 i_1085 (.A(n_1991), .ZN(n_1990));
   OAI21_X1 i_1086 (.A(n_2258), .B1(n_2203), .B2(n_1992), .ZN(n_1991));
   AOI21_X1 i_1087 (.A(n_2262), .B1(n_2205), .B2(n_2014), .ZN(n_1992));
   OAI21_X1 i_1088 (.A(n_2205), .B1(n_379), .B2(n_418), .ZN(n_1993));
   AOI21_X1 i_1089 (.A(n_2261), .B1(n_505), .B2(n_550), .ZN(n_1994));
   XOR2_X1 i_1090 (.A(n_2012), .B(n_2001), .Z(out31[25]));
   XOR2_X1 i_1091 (.A(n_2000), .B(n_1997), .Z(out31[26]));
   XOR2_X1 i_1092 (.A(n_1998), .B(n_1995), .Z(out31[27]));
   NOR2_X1 i_1093 (.A1(n_2240), .A2(n_2213), .ZN(n_1995));
   XNOR2_X1 i_1094 (.A(n_2002), .B(n_1996), .ZN(out31[28]));
   OAI21_X1 i_1095 (.A(n_2239), .B1(n_2213), .B2(n_1998), .ZN(n_1996));
   NOR2_X1 i_1096 (.A1(n_2242), .A2(n_2215), .ZN(n_1997));
   INV_X1 i_1097 (.A(n_1999), .ZN(n_1998));
   OAI21_X1 i_1098 (.A(n_2241), .B1(n_2215), .B2(n_2000), .ZN(n_1999));
   AOI21_X1 i_1099 (.A(n_2237), .B1(n_2217), .B2(n_2012), .ZN(n_2000));
   OAI21_X1 i_1100 (.A(n_2217), .B1(n_596), .B2(n_598), .ZN(n_2001));
   AOI21_X1 i_1101 (.A(n_2244), .B1(n_701), .B2(n_754), .ZN(n_2002));
   XOR2_X1 i_1102 (.A(n_2010), .B(n_2009), .Z(out31[29]));
   XOR2_X1 i_1103 (.A(n_2008), .B(n_2005), .Z(out31[30]));
   XOR2_X1 i_1104 (.A(n_2006), .B(n_2003), .Z(out31[31]));
   NOR2_X1 i_1105 (.A1(n_2249), .A2(n_2207), .ZN(n_2003));
   XOR2_X1 i_1106 (.A(n_2016), .B(n_2004), .Z(out31[32]));
   OAI21_X1 i_1107 (.A(n_2248), .B1(n_2207), .B2(n_2006), .ZN(n_2004));
   NOR2_X1 i_1108 (.A1(n_2251), .A2(n_2210), .ZN(n_2005));
   INV_X1 i_1109 (.A(n_2007), .ZN(n_2006));
   OAI21_X1 i_1110 (.A(n_2250), .B1(n_2210), .B2(n_2008), .ZN(n_2007));
   AOI21_X1 i_1111 (.A(n_2246), .B1(n_2211), .B2(n_2010), .ZN(n_2008));
   OAI21_X1 i_1112 (.A(n_2211), .B1(n_755), .B2(n_810), .ZN(n_2009));
   INV_X1 i_1113 (.A(n_2011), .ZN(n_2010));
   OAI21_X1 i_1114 (.A(n_2212), .B1(n_2236), .B2(n_2012), .ZN(n_2011));
   INV_X1 i_1115 (.A(n_2013), .ZN(n_2012));
   OAI21_X1 i_1116 (.A(n_2200), .B1(n_2254), .B2(n_2014), .ZN(n_2013));
   INV_X1 i_1117 (.A(n_2015), .ZN(n_2014));
   OAI21_X1 i_1118 (.A(n_2218), .B1(n_2263), .B2(n_2225), .ZN(n_2015));
   OAI21_X1 i_1119 (.A(n_2252), .B1(n_2328), .B2(n_2327), .ZN(n_2016));
   XOR2_X1 i_1120 (.A(n_2198), .B(n_2023), .Z(out31[33]));
   XOR2_X1 i_1121 (.A(n_2022), .B(n_2019), .Z(out31[34]));
   XOR2_X1 i_1122 (.A(n_2020), .B(n_2017), .Z(out31[35]));
   NOR2_X1 i_1123 (.A1(n_2167), .A2(n_2157), .ZN(n_2017));
   XNOR2_X1 i_1124 (.A(n_2024), .B(n_2018), .ZN(out31[36]));
   OAI21_X1 i_1125 (.A(n_2166), .B1(n_2157), .B2(n_2020), .ZN(n_2018));
   NOR2_X1 i_1126 (.A1(n_2169), .A2(n_2159), .ZN(n_2019));
   INV_X1 i_1127 (.A(n_2021), .ZN(n_2020));
   OAI21_X1 i_1128 (.A(n_2168), .B1(n_2159), .B2(n_2022), .ZN(n_2021));
   AOI21_X1 i_1129 (.A(n_2164), .B1(n_2198), .B2(n_2161), .ZN(n_2022));
   OAI21_X1 i_1130 (.A(n_2161), .B1(n_987), .B2(n_1044), .ZN(n_2023));
   AOI21_X1 i_1131 (.A(n_2171), .B1(n_1155), .B2(n_1206), .ZN(n_2024));
   XOR2_X1 i_1132 (.A(n_2052), .B(n_2031), .Z(out31[37]));
   OAI21_X1 i_1142 (.A(n_2154), .B1(n_1207), .B2(n_1256), .ZN(n_2031));
   XOR2_X1 i_1144 (.A(n_2050), .B(n_2039), .Z(out31[41]));
   OAI21_X1 i_1154 (.A(n_2140), .B1(n_1395), .B2(n_1436), .ZN(n_2039));
   XOR2_X1 i_1174 (.A(n_2133), .B(n_2061), .Z(out31[49]));
   XOR2_X1 i_1175 (.A(n_2060), .B(n_2057), .Z(out31[50]));
   AOI21_X1 i_1180 (.A(n_2131), .B1(n_1701), .B2(n_1724), .ZN(n_2057));
   OAI21_X1 i_1184 (.A(n_2126), .B1(n_1675), .B2(n_1700), .ZN(n_2061));
   XOR2_X1 i_1186 (.A(n_2119), .B(n_2069), .Z(out31[53]));
   OAI21_X1 i_1196 (.A(n_2102), .B1(n_1767), .B2(n_1784), .ZN(n_2069));
   XNOR2_X1 i_1198 (.A(n_2079), .B(n_2078), .ZN(out31[57]));
   OAI21_X1 i_1209 (.A(n_2095), .B1(n_1827), .B2(n_1836), .ZN(n_2078));
   OAI21_X1 i_1226 (.A(n_2114), .B1(n_2094), .B2(n_2093), .ZN(n_2092));
   AOI21_X1 i_1233 (.A(n_2106), .B1(n_2102), .B2(n_2101), .ZN(n_2099));
   NAND3_X1 i_1240 (.A1(n_2111), .A2(n_2107), .A3(n_2109), .ZN(n_2106));
   INV_X1 i_1245 (.A(n_2112), .ZN(n_2111));
   NOR2_X1 i_1246 (.A1(n_1815), .A2(n_1826), .ZN(n_2112));
   NOR3_X1 i_1248 (.A1(n_2118), .A2(n_2116), .A3(n_2117), .ZN(n_2114));
   NOR2_X1 i_1250 (.A1(n_1845), .A2(n_1850), .ZN(n_2116));
   NOR2_X1 i_1251 (.A1(n_1837), .A2(n_1844), .ZN(n_2117));
   NOR2_X1 i_1252 (.A1(n_1851), .A2(n_1854), .ZN(n_2118));
   NOR2_X1 i_1264 (.A1(n_1725), .A2(n_1746), .ZN(n_2130));
   NOR2_X1 i_1266 (.A1(n_1747), .A2(n_1766), .ZN(n_2132));
   OAI21_X1 i_1276 (.A(n_2145), .B1(n_2188), .B2(n_2144), .ZN(n_2142));
   OAI21_X1 i_1279 (.A(n_2184), .B1(n_2147), .B2(n_2146), .ZN(n_2145));
   INV_X1 i_1293 (.A(n_2160), .ZN(n_2159));
   NOR2_X1 i_1298 (.A1(n_987), .A2(n_1044), .ZN(n_2164));
   NOR3_X1 i_1318 (.A1(n_2188), .A2(n_2186), .A3(n_2187), .ZN(n_2184));
   NOR2_X1 i_1320 (.A1(n_1617), .A2(n_1646), .ZN(n_2186));
   NOR2_X1 i_1321 (.A1(n_1585), .A2(n_1616), .ZN(n_2187));
   NOR2_X1 i_1322 (.A1(n_1647), .A2(n_1674), .ZN(n_2188));
   AND2_X1 i_1335 (.A1(n_461), .A2(n_504), .ZN(n_2201));
   AOI21_X1 i_1336 (.A(n_2255), .B1(n_2205), .B2(n_2204), .ZN(n_2202));
   INV_X1 i_1337 (.A(n_2204), .ZN(n_2203));
   NAND2_X1 i_1338 (.A1(n_419), .A2(n_460), .ZN(n_2204));
   NAND2_X1 i_1339 (.A1(n_379), .A2(n_418), .ZN(n_2205));
   INV_X1 i_1341 (.A(n_2208), .ZN(n_2207));
   AND2_X1 i_1344 (.A1(n_811), .A2(n_868), .ZN(n_2210));
   NAND2_X1 i_1345 (.A1(n_755), .A2(n_810), .ZN(n_2211));
   INV_X1 i_1349 (.A(n_2216), .ZN(n_2215));
   AND2_X1 i_1353 (.A1(n_305), .A2(n_340), .ZN(n_2219));
   INV_X1 i_1355 (.A(n_2222), .ZN(n_2221));
   NOR2_X1 i_1360 (.A1(n_268), .A2(n_270), .ZN(n_2226));
   NOR2_X1 i_1363 (.A1(n_305), .A2(n_340), .ZN(n_2229));
   NOR2_X1 i_1365 (.A1(n_271), .A2(n_304), .ZN(n_2231));
   NOR2_X1 i_1371 (.A1(n_596), .A2(n_598), .ZN(n_2237));
   NOR2_X1 i_1374 (.A1(n_649), .A2(n_700), .ZN(n_2240));
   NOR2_X1 i_1376 (.A1(n_599), .A2(n_648), .ZN(n_2242));
   NAND3_X1 i_1389 (.A1(n_2260), .A2(n_2256), .A3(n_2258), .ZN(n_2255));
   INV_X1 i_1390 (.A(n_2257), .ZN(n_2256));
   NOR2_X1 i_1391 (.A1(n_461), .A2(n_504), .ZN(n_2257));
   INV_X1 i_1392 (.A(n_2259), .ZN(n_2258));
   NOR2_X1 i_1393 (.A1(n_419), .A2(n_460), .ZN(n_2259));
   INV_X1 i_1394 (.A(n_2261), .ZN(n_2260));
   NOR2_X1 i_1395 (.A1(n_505), .A2(n_550), .ZN(n_2261));
   NOR2_X1 i_1396 (.A1(n_379), .A2(n_418), .ZN(n_2262));
   NOR2_X1 i_1398 (.A1(n_2276), .A2(n_2266), .ZN(n_2264));
   INV_X1 i_1399 (.A(n_2266), .ZN(n_2265));
   NAND2_X1 i_1400 (.A1(n_206), .A2(n_208), .ZN(n_2266));
   AND2_X1 i_1401 (.A1(n_236), .A2(n_238), .ZN(n_2267));
   AOI21_X1 i_1402 (.A(n_2273), .B1(n_2270), .B2(n_2269), .ZN(n_2268));
   NAND2_X1 i_1403 (.A1(n_178), .A2(n_180), .ZN(n_2269));
   NAND2_X1 i_1404 (.A1(n_152), .A2(n_154), .ZN(n_2270));
   NOR3_X1 i_1405 (.A1(n_2273), .A2(n_2272), .A3(n_2277), .ZN(n_2271));
   NOR2_X1 i_1406 (.A1(n_152), .A2(n_154), .ZN(n_2272));
   OR3_X1 i_1407 (.A1(n_2276), .A2(n_2274), .A3(n_2275), .ZN(n_2273));
   NOR2_X1 i_1408 (.A1(n_206), .A2(n_208), .ZN(n_2274));
   NOR2_X1 i_1409 (.A1(n_178), .A2(n_180), .ZN(n_2275));
   NOR2_X1 i_1410 (.A1(n_236), .A2(n_238), .ZN(n_2276));
   NOR4_X1 i_1411 (.A1(n_2281), .A2(n_2278), .A3(n_2282), .A4(n_2285), .ZN(
      n_2277));
   NOR2_X1 i_1412 (.A1(n_2290), .A2(n_2280), .ZN(n_2278));
   INV_X1 i_1413 (.A(n_2280), .ZN(n_2279));
   NAND2_X1 i_1414 (.A1(n_106), .A2(n_108), .ZN(n_2280));
   AND2_X1 i_1415 (.A1(n_128), .A2(n_130), .ZN(n_2281));
   AOI21_X1 i_1416 (.A(n_2287), .B1(n_2284), .B2(n_2283), .ZN(n_2282));
   NAND2_X1 i_1417 (.A1(n_86), .A2(n_88), .ZN(n_2283));
   NAND2_X1 i_1418 (.A1(n_68), .A2(n_70), .ZN(n_2284));
   NOR3_X1 i_1419 (.A1(n_2287), .A2(n_2286), .A3(n_2291), .ZN(n_2285));
   NOR2_X1 i_1420 (.A1(n_68), .A2(n_70), .ZN(n_2286));
   OR3_X1 i_1421 (.A1(n_2290), .A2(n_2288), .A3(n_2289), .ZN(n_2287));
   NOR2_X1 i_1422 (.A1(n_106), .A2(n_108), .ZN(n_2288));
   NOR2_X1 i_1423 (.A1(n_86), .A2(n_88), .ZN(n_2289));
   NOR2_X1 i_1424 (.A1(n_128), .A2(n_130), .ZN(n_2290));
   NOR4_X1 i_1425 (.A1(n_2295), .A2(n_2292), .A3(n_2296), .A4(n_2299), .ZN(
      n_2291));
   NOR2_X1 i_1426 (.A1(n_2304), .A2(n_2294), .ZN(n_2292));
   INV_X1 i_1427 (.A(n_2294), .ZN(n_2293));
   NAND2_X1 i_1428 (.A1(n_38), .A2(n_40), .ZN(n_2294));
   AND2_X1 i_1429 (.A1(n_52), .A2(n_54), .ZN(n_2295));
   AOI21_X1 i_1430 (.A(n_2301), .B1(n_2298), .B2(n_2297), .ZN(n_2296));
   NAND2_X1 i_1431 (.A1(n_26), .A2(n_28), .ZN(n_2297));
   NAND2_X1 i_1432 (.A1(n_16), .A2(n_18), .ZN(n_2298));
   NOR3_X1 i_1433 (.A1(n_2301), .A2(n_2300), .A3(n_2305), .ZN(n_2299));
   NOR2_X1 i_1434 (.A1(n_16), .A2(n_18), .ZN(n_2300));
   OR3_X1 i_1435 (.A1(n_2304), .A2(n_2302), .A3(n_2303), .ZN(n_2301));
   NOR2_X1 i_1436 (.A1(n_38), .A2(n_40), .ZN(n_2302));
   NOR2_X1 i_1437 (.A1(n_26), .A2(n_28), .ZN(n_2303));
   NOR2_X1 i_1438 (.A1(n_52), .A2(n_54), .ZN(n_2304));
   NAND2_X1 i_1439 (.A1(n_2314), .A2(n_2306), .ZN(n_2305));
   OAI21_X1 i_1440 (.A(n_2307), .B1(n_2330), .B2(n_2329), .ZN(n_2306));
   OAI22_X1 i_1441 (.A1(n_2), .A2(n_4), .B1(n_2312), .B2(n_2308), .ZN(n_2307));
   AOI21_X1 i_1442 (.A(n_2311), .B1(n_2310), .B2(n_2309), .ZN(n_2308));
   NAND2_X1 i_1443 (.A1(out[2]), .A2(n_0), .ZN(n_2309));
   NAND2_X1 i_1444 (.A1(p_0[1]), .A2(out[1]), .ZN(n_2310));
   NOR2_X1 i_1445 (.A1(out[2]), .A2(n_0), .ZN(n_2311));
   INV_X1 i_1446 (.A(n_2313), .ZN(n_2312));
   NAND2_X1 i_1447 (.A1(n_2), .A2(n_4), .ZN(n_2313));
   NAND2_X1 i_1448 (.A1(n_2330), .A2(n_2329), .ZN(n_2314));
   OR3_X1 i_1451 (.A1(n_2331), .A2(n_2320), .A3(p_29[62]), .ZN(n_2317));
   OAI22_X1 i_1452 (.A1(n_2331), .A2(n_2320), .B1(p_29[62]), .B2(n_2319), 
      .ZN(n_2318));
   AND2_X1 i_1453 (.A1(n_2331), .A2(n_2320), .ZN(n_2319));
   OAI22_X1 i_1454 (.A1(p_29[61]), .A2(n_2321), .B1(n_2335), .B2(p_30[61]), 
      .ZN(n_2320));
   INV_X1 i_1455 (.A(n_2322), .ZN(n_2321));
   NAND2_X1 i_1456 (.A1(n_2335), .A2(p_30[61]), .ZN(n_2322));
   INV_X1 i_1458 (.A(n_1854), .ZN(n_2324));
   INV_X1 i_1460 (.A(n_1851), .ZN(n_2326));
   INV_X1 i_1462 (.A(n_929), .ZN(n_2328));
   INV_X1 i_1463 (.A(n_10), .ZN(n_2329));
   INV_X1 i_1464 (.A(n_6), .ZN(n_2330));
   INV_X1 i_1465 (.A(p_30[62]), .ZN(n_2331));
   INV_X1 i_1466 (.A(p_29[60]), .ZN(n_2332));
   INV_X1 i_1467 (.A(p_28[59]), .ZN(n_2333));
   INV_X1 i_1468 (.A(p_28[60]), .ZN(n_2334));
   INV_X1 i_1469 (.A(p_28[61]), .ZN(n_2335));
   INV_X1 i_1470 (.A(p_27[58]), .ZN(n_2336));
   INV_X1 i_1471 (.A(p_27[59]), .ZN(n_2337));
   INV_X1 i_1472 (.A(p_26[57]), .ZN(n_2338));
   INV_X1 i_1473 (.A(p_26[58]), .ZN(n_2339));
   INV_X1 i_1474 (.A(p_25[56]), .ZN(n_2340));
   INV_X1 i_1475 (.A(p_25[57]), .ZN(n_2341));
   INV_X1 i_1476 (.A(p_24[55]), .ZN(n_2342));
   INV_X1 i_1477 (.A(p_24[56]), .ZN(n_2343));
   INV_X1 i_1478 (.A(p_23[54]), .ZN(n_2344));
   INV_X1 i_1479 (.A(p_23[55]), .ZN(n_2345));
   INV_X1 i_1480 (.A(p_22[53]), .ZN(n_2346));
   INV_X1 i_1481 (.A(p_22[54]), .ZN(n_2347));
   INV_X1 i_1482 (.A(p_21[52]), .ZN(n_2348));
   INV_X1 i_1483 (.A(p_21[53]), .ZN(n_2349));
   INV_X1 i_1484 (.A(p_20[51]), .ZN(n_2350));
   INV_X1 i_1485 (.A(p_20[52]), .ZN(n_2351));
   INV_X1 i_1486 (.A(p_19[50]), .ZN(n_2352));
   INV_X1 i_1487 (.A(p_19[51]), .ZN(n_2353));
   INV_X1 i_1488 (.A(p_18[49]), .ZN(n_2354));
   INV_X1 i_1489 (.A(p_18[50]), .ZN(n_2355));
   INV_X1 i_1490 (.A(p_17[48]), .ZN(n_2356));
   INV_X1 i_1491 (.A(p_17[49]), .ZN(n_2357));
   INV_X1 i_1492 (.A(p_16[47]), .ZN(n_2358));
   INV_X1 i_1493 (.A(p_16[48]), .ZN(n_2359));
   INV_X1 i_1494 (.A(p_15[46]), .ZN(n_2360));
   INV_X1 i_1495 (.A(p_15[47]), .ZN(n_2361));
   INV_X1 i_1496 (.A(p_14[45]), .ZN(n_2362));
   INV_X1 i_1497 (.A(p_14[46]), .ZN(n_2363));
   INV_X1 i_1498 (.A(p_13[44]), .ZN(n_2364));
   INV_X1 i_1499 (.A(p_13[45]), .ZN(n_2365));
   INV_X1 i_1500 (.A(p_12[43]), .ZN(n_2366));
   INV_X1 i_1501 (.A(p_12[44]), .ZN(n_2367));
   INV_X1 i_1502 (.A(p_11[42]), .ZN(n_2368));
   INV_X1 i_1503 (.A(p_11[43]), .ZN(n_2369));
   INV_X1 i_1504 (.A(p_10[41]), .ZN(n_2370));
   INV_X1 i_1505 (.A(p_10[42]), .ZN(n_2371));
   INV_X1 i_1506 (.A(p_9[40]), .ZN(n_2372));
   INV_X1 i_1507 (.A(p_9[41]), .ZN(n_2373));
   INV_X1 i_1509 (.A(p_8[40]), .ZN(n_2375));
   INV_X1 i_1516 (.A(p_4[35]), .ZN(n_2382));
   INV_X1 i_1519 (.A(p_3[35]), .ZN(n_2385));
   INV_X1 i_1522 (.A(p_1[32]), .ZN(n_2388));
   INV_X1 i_1523 (.A(p_1[33]), .ZN(n_2389));
   INV_X1 i_1524 (.A(p_0[32]), .ZN(n_2390));
   INV_X1 i_994 (.A(n_1856), .ZN(n_2323));
   INV_X1 i_995 (.A(n_1855), .ZN(n_2325));
   INV_X1 i_996 (.A(n_2026), .ZN(n_2123));
   NAND2_X1 i_999 (.A1(n_2040), .A2(n_2041), .ZN(n_2225));
   INV_X1 i_1000 (.A(n_2055), .ZN(n_2218));
   NAND2_X1 i_1001 (.A1(n_2045), .A2(n_2044), .ZN(n_2254));
   INV_X1 i_1002 (.A(n_2499), .ZN(n_2212));
   INV_X1 i_1005 (.A(n_2251), .ZN(n_2250));
   INV_X1 i_1009 (.A(n_2249), .ZN(n_2248));
   INV_X1 i_1010 (.A(n_2113), .ZN(n_2213));
   INV_X1 i_1011 (.A(n_2034), .ZN(n_2263));
   OAI221_X1 i_1012 (.A(n_2092), .B1(n_2090), .B2(n_2118), .C1(n_2326), .C2(
      n_2324), .ZN(n_1924));
   INV_X1 i_1013 (.A(n_2097), .ZN(n_1930));
   INV_X1 i_1017 (.A(n_1942), .ZN(n_1939));
   OAI21_X1 i_1018 (.A(n_2114), .B1(n_1827), .B2(n_1836), .ZN(n_1942));
   INV_X1 i_1019 (.A(n_2106), .ZN(n_1948));
   INV_X1 i_1133 (.A(n_2105), .ZN(n_2025));
   NAND2_X1 i_1134 (.A1(n_1747), .A2(n_1766), .ZN(n_2026));
   NAND2_X1 i_1135 (.A1(n_2029), .A2(n_2028), .ZN(n_2027));
   NAND2_X1 i_1136 (.A1(n_2125), .A2(n_2126), .ZN(n_2028));
   NOR3_X1 i_1137 (.A1(n_2131), .A2(n_2130), .A3(n_2132), .ZN(n_2029));
   NAND2_X1 i_1138 (.A1(n_648), .A2(n_599), .ZN(n_2216));
   NAND2_X1 i_1139 (.A1(n_598), .A2(n_596), .ZN(n_2217));
   AND2_X1 i_1140 (.A1(n_2032), .A2(n_2030), .ZN(n_2200));
   AOI22_X1 i_1141 (.A1(n_2260), .A2(n_2201), .B1(n_505), .B2(n_550), .ZN(n_2030));
   INV_X1 i_1143 (.A(n_2202), .ZN(n_2032));
   NAND3_X1 i_1145 (.A1(n_2040), .A2(n_2041), .A3(n_2034), .ZN(n_2033));
   NAND4_X1 i_1146 (.A1(n_2036), .A2(n_2035), .A3(n_2038), .A4(n_2037), .ZN(
      n_2034));
   INV_X1 i_1147 (.A(n_2271), .ZN(n_2035));
   INV_X1 i_1148 (.A(n_2268), .ZN(n_2036));
   INV_X1 i_1149 (.A(n_2264), .ZN(n_2037));
   INV_X1 i_1150 (.A(n_2267), .ZN(n_2038));
   INV_X1 i_1151 (.A(n_2227), .ZN(n_2040));
   INV_X1 i_1152 (.A(n_2226), .ZN(n_2041));
   NAND4_X1 i_1153 (.A1(n_2104), .A2(n_2239), .A3(n_2241), .A4(n_2042), .ZN(
      n_2236));
   INV_X1 i_1155 (.A(n_2237), .ZN(n_2042));
   AOI22_X1 i_1156 (.A1(n_2318), .A2(n_2317), .B1(p_29[62]), .B2(n_2319), 
      .ZN(n_2043));
   INV_X1 i_1157 (.A(n_2262), .ZN(n_2044));
   INV_X1 i_1158 (.A(n_2255), .ZN(n_2045));
   INV_X1 i_1159 (.A(n_2095), .ZN(n_2094));
   OAI21_X1 i_1160 (.A(n_2097), .B1(n_2119), .B2(n_2085), .ZN(n_2079));
   INV_X1 i_1161 (.A(n_2101), .ZN(n_2100));
   INV_X1 i_1162 (.A(n_2122), .ZN(n_2121));
   INV_X1 i_1163 (.A(n_2062), .ZN(n_2060));
   INV_X1 i_1164 (.A(n_2148), .ZN(n_2147));
   INV_X1 i_1165 (.A(n_2139), .ZN(n_2138));
   INV_X1 i_1166 (.A(n_2463), .ZN(n_2157));
   INV_X1 i_1167 (.A(n_2144), .ZN(n_2046));
   NAND2_X1 i_1168 (.A1(n_1674), .A2(n_1647), .ZN(n_2047));
   INV_X1 i_1169 (.A(n_2188), .ZN(n_2048));
   INV_X1 i_1170 (.A(n_1844), .ZN(n_2049));
   INV_X1 i_1171 (.A(n_1837), .ZN(n_2051));
   OR2_X1 i_1172 (.A1(n_2093), .A2(n_2117), .ZN(n_2053));
   INV_X1 i_1173 (.A(n_2055), .ZN(n_2054));
   OAI21_X1 i_1176 (.A(n_2058), .B1(n_2233), .B2(n_2056), .ZN(n_2055));
   AOI21_X1 i_1177 (.A(n_2219), .B1(n_378), .B2(n_376), .ZN(n_2056));
   OR2_X1 i_1178 (.A1(n_2227), .A2(n_2059), .ZN(n_2058));
   AND2_X1 i_1179 (.A1(n_2222), .A2(n_2223), .ZN(n_2059));
   NAND2_X1 i_1181 (.A1(n_304), .A2(n_271), .ZN(n_2222));
   NAND2_X1 i_1182 (.A1(n_270), .A2(n_268), .ZN(n_2223));
   OAI211_X1 i_1183 (.A(n_2228), .B(n_2230), .C1(n_378), .C2(n_376), .ZN(n_2227));
   INV_X1 i_1185 (.A(n_2231), .ZN(n_2230));
   INV_X1 i_1187 (.A(n_2229), .ZN(n_2228));
   NOR2_X1 i_1188 (.A1(n_378), .A2(n_376), .ZN(n_2233));
   INV_X1 i_1189 (.A(n_2316), .ZN(n_2062));
   INV_X1 i_1190 (.A(n_2110), .ZN(n_2109));
   INV_X1 i_1191 (.A(n_2406), .ZN(n_2093));
   INV_X1 i_1192 (.A(n_2206), .ZN(n_2050));
   INV_X1 i_1193 (.A(n_2169), .ZN(n_2168));
   INV_X1 i_1194 (.A(n_2167), .ZN(n_2166));
   INV_X1 i_1195 (.A(n_2484), .ZN(n_2198));
   XNOR2_X1 i_1197 (.A(n_2063), .B(p_8[39]), .ZN(n_1923));
   XNOR2_X1 i_1199 (.A(n_2120), .B(p_7[39]), .ZN(n_2063));
   XNOR2_X1 i_1200 (.A(n_2064), .B(p_6[37]), .ZN(n_1929));
   XNOR2_X1 i_1201 (.A(n_2103), .B(p_4[59]), .ZN(n_2064));
   INV_X1 i_1202 (.A(n_2065), .ZN(out31[38]));
   XOR2_X1 i_1203 (.A(n_2066), .B(n_2071), .Z(n_2065));
   NAND2_X1 i_1204 (.A1(n_2153), .A2(n_2072), .ZN(n_2066));
   XOR2_X1 i_1205 (.A(n_2067), .B(n_2070), .Z(out31[39]));
   NAND2_X1 i_1206 (.A1(n_2108), .A2(n_2191), .ZN(n_2067));
   XNOR2_X1 i_1207 (.A(n_2068), .B(n_2074), .ZN(out31[40]));
   AOI22_X1 i_1208 (.A1(n_2070), .A2(n_2108), .B1(n_2483), .B2(n_2482), .ZN(
      n_2068));
   OAI21_X1 i_1210 (.A(n_2072), .B1(n_2071), .B2(n_2073), .ZN(n_2070));
   OAI21_X1 i_1211 (.A(n_2154), .B1(n_2052), .B2(n_2098), .ZN(n_2071));
   INV_X1 i_1212 (.A(n_2096), .ZN(n_2072));
   INV_X1 i_1213 (.A(n_2153), .ZN(n_2073));
   XNOR2_X1 i_1214 (.A(n_1394), .B(n_1351), .ZN(n_2074));
   XNOR2_X1 i_1215 (.A(n_2091), .B(n_2075), .ZN(out31[42]));
   NOR2_X1 i_1216 (.A1(n_2138), .A2(n_2474), .ZN(n_2075));
   XOR2_X1 i_1217 (.A(n_2076), .B(n_2199), .Z(out31[45]));
   NAND2_X1 i_1218 (.A1(n_2077), .A2(n_2148), .ZN(n_2076));
   INV_X1 i_1219 (.A(n_2232), .ZN(n_2077));
   INV_X1 i_1220 (.A(n_2224), .ZN(n_2146));
   NAND2_X1 i_1221 (.A1(n_2048), .A2(n_2047), .ZN(n_2080));
   XNOR2_X1 i_1222 (.A(n_2247), .B(n_2081), .ZN(out31[51]));
   NOR2_X1 i_1223 (.A1(n_2121), .A2(n_2130), .ZN(n_2081));
   NOR2_X1 i_1224 (.A1(n_1724), .A2(n_1701), .ZN(n_2131));
   NAND2_X1 i_1225 (.A1(n_1724), .A2(n_1701), .ZN(n_2125));
   XNOR2_X1 i_1227 (.A(n_2396), .B(n_2082), .ZN(out31[54]));
   NOR2_X1 i_1228 (.A1(n_2110), .A2(n_2100), .ZN(n_2082));
   NOR2_X1 i_1229 (.A1(n_1784), .A2(n_1767), .ZN(n_2105));
   NAND2_X1 i_1230 (.A1(n_1784), .A2(n_1767), .ZN(n_2102));
   OR2_X1 i_1231 (.A1(n_1827), .A2(n_1836), .ZN(n_2083));
   AOI221_X1 i_1232 (.A(n_2099), .B1(n_1815), .B2(n_1826), .C1(n_2111), .C2(
      n_2400), .ZN(n_2097));
   NAND2_X1 i_1234 (.A1(n_1814), .A2(n_1801), .ZN(n_2084));
   NAND2_X1 i_1235 (.A1(n_1827), .A2(n_1836), .ZN(n_2095));
   NAND2_X1 i_1236 (.A1(n_1948), .A2(n_2025), .ZN(n_2085));
   NAND2_X1 i_1237 (.A1(n_2323), .A2(n_2325), .ZN(n_2086));
   NAND2_X1 i_1238 (.A1(n_2508), .A2(n_2509), .ZN(n_2087));
   OAI211_X1 i_1239 (.A(n_2027), .B(n_2026), .C1(n_2132), .C2(n_2122), .ZN(
      n_2088));
   NAND2_X1 i_1241 (.A1(n_1856), .A2(n_1855), .ZN(n_2089));
   NOR2_X1 i_1242 (.A1(n_2173), .A2(n_2175), .ZN(n_2091));
   NOR2_X1 i_1243 (.A1(n_1304), .A2(n_1257), .ZN(n_2096));
   NOR2_X1 i_1244 (.A1(n_1256), .A2(n_1207), .ZN(n_2098));
   INV_X1 i_1247 (.A(p_5[37]), .ZN(n_2103));
   INV_X1 i_1249 (.A(n_2244), .ZN(n_2104));
   NAND2_X1 i_1253 (.A1(n_1350), .A2(n_1305), .ZN(n_2108));
   NAND2_X1 i_1254 (.A1(n_700), .A2(n_649), .ZN(n_2113));
   NAND2_X1 i_1255 (.A1(n_2482), .A2(n_2483), .ZN(n_2191));
   INV_X1 i_1256 (.A(n_2439), .ZN(n_2119));
   OAI21_X1 i_1257 (.A(n_2115), .B1(p_6[59]), .B2(n_2124), .ZN(n_1925));
   OAI21_X1 i_1258 (.A(p_7[39]), .B1(n_2120), .B2(p_8[39]), .ZN(n_2115));
   INV_X1 i_1259 (.A(p_6[59]), .ZN(n_2120));
   INV_X1 i_1260 (.A(p_8[39]), .ZN(n_2124));
   OAI21_X1 i_1261 (.A(n_2127), .B1(p_5[59]), .B2(n_2376), .ZN(n_1928));
   OAI21_X1 i_1262 (.A(p_6[38]), .B1(n_2128), .B2(p_7[38]), .ZN(n_2127));
   INV_X1 i_1263 (.A(p_5[59]), .ZN(n_2128));
   INV_X1 i_1265 (.A(p_7[38]), .ZN(n_2376));
   AOI21_X1 i_1267 (.A(n_2129), .B1(p_4[59]), .B2(n_2134), .ZN(n_1931));
   NOR2_X1 i_1268 (.A1(p_5[37]), .A2(p_6[37]), .ZN(n_2129));
   NAND2_X1 i_1269 (.A1(p_5[37]), .A2(p_6[37]), .ZN(n_2134));
   OAI21_X1 i_1270 (.A(n_2135), .B1(p_3[59]), .B2(n_2380), .ZN(n_1934));
   OAI21_X1 i_1271 (.A(p_4[36]), .B1(n_2136), .B2(p_5[36]), .ZN(n_2135));
   INV_X1 i_1272 (.A(p_3[59]), .ZN(n_2136));
   INV_X1 i_1273 (.A(p_5[36]), .ZN(n_2380));
   NAND2_X1 i_1274 (.A1(n_2149), .A2(n_2137), .ZN(n_1940));
   NAND2_X1 i_1275 (.A1(n_2143), .A2(p_3[34]), .ZN(n_2137));
   XNOR2_X1 i_1277 (.A(n_2141), .B(p_3[34]), .ZN(n_1938));
   NAND2_X1 i_1278 (.A1(n_2149), .A2(n_2143), .ZN(n_2141));
   NAND2_X1 i_1280 (.A1(p_1[59]), .A2(n_2150), .ZN(n_2143));
   OR2_X1 i_1281 (.A1(p_1[59]), .A2(n_2150), .ZN(n_2149));
   INV_X1 i_1282 (.A(p_2[34]), .ZN(n_2150));
   XNOR2_X1 i_1283 (.A(n_2151), .B(p_0[59]), .ZN(n_1941));
   XNOR2_X1 i_1284 (.A(n_2386), .B(p_1[33]), .ZN(n_2151));
   INV_X1 i_1285 (.A(p_2[33]), .ZN(n_2386));
   OAI21_X1 i_1286 (.A(n_1947), .B1(out[61]), .B2(n_2152), .ZN(n_1946));
   NOR2_X1 i_1287 (.A1(p_29[32]), .A2(p_30[32]), .ZN(n_2152));
   NAND2_X1 i_1288 (.A1(p_29[32]), .A2(p_30[32]), .ZN(n_1947));
   XNOR2_X1 i_1289 (.A(n_2156), .B(n_2155), .ZN(out31[43]));
   NAND2_X1 i_1290 (.A1(n_2179), .A2(n_2448), .ZN(n_2155));
   NAND2_X1 i_1291 (.A1(n_2172), .A2(n_2139), .ZN(n_2156));
   NAND2_X1 i_1292 (.A1(n_2158), .A2(n_2165), .ZN(out31[44]));
   OAI21_X1 i_1294 (.A(n_2163), .B1(n_2162), .B2(n_2475), .ZN(n_2158));
   INV_X1 i_1295 (.A(n_2170), .ZN(n_2162));
   INV_X1 i_1296 (.A(n_2177), .ZN(n_2163));
   NAND3_X1 i_1297 (.A1(n_2170), .A2(n_2179), .A3(n_2177), .ZN(n_2165));
   NAND3_X1 i_1299 (.A1(n_2172), .A2(n_2139), .A3(n_2448), .ZN(n_2170));
   OAI21_X1 i_1300 (.A(n_2176), .B1(n_2173), .B2(n_2175), .ZN(n_2172));
   INV_X1 i_1301 (.A(n_2174), .ZN(n_2173));
   NAND2_X1 i_1302 (.A1(n_2206), .A2(n_2476), .ZN(n_2174));
   INV_X1 i_1303 (.A(n_2140), .ZN(n_2175));
   INV_X1 i_1304 (.A(n_2474), .ZN(n_2176));
   NAND2_X1 i_1305 (.A1(n_2178), .A2(n_2449), .ZN(n_2177));
   INV_X1 i_1306 (.A(n_2473), .ZN(n_2178));
   INV_X1 i_1307 (.A(n_2475), .ZN(n_2179));
   XNOR2_X1 i_1308 (.A(n_2181), .B(n_2180), .ZN(out31[46]));
   OR2_X1 i_1309 (.A1(n_2146), .A2(n_2187), .ZN(n_2180));
   OAI21_X1 i_1310 (.A(n_2148), .B1(n_2199), .B2(n_2232), .ZN(n_2181));
   NAND2_X1 i_1311 (.A1(n_2182), .A2(n_2185), .ZN(out31[47]));
   NAND2_X1 i_1312 (.A1(n_2183), .A2(n_2190), .ZN(n_2182));
   OAI21_X1 i_1313 (.A(n_2197), .B1(n_1585), .B2(n_1616), .ZN(n_2183));
   OAI211_X1 i_1314 (.A(n_2197), .B(n_2189), .C1(n_1585), .C2(n_1616), .ZN(
      n_2185));
   INV_X1 i_1315 (.A(n_2190), .ZN(n_2189));
   NOR2_X1 i_1316 (.A1(n_2186), .A2(n_2046), .ZN(n_2190));
   NAND2_X1 i_1317 (.A1(n_2192), .A2(n_2194), .ZN(out31[48]));
   NAND2_X1 i_1319 (.A1(n_2193), .A2(n_2080), .ZN(n_2192));
   NAND2_X1 i_1323 (.A1(n_2195), .A2(n_2144), .ZN(n_2193));
   NAND3_X1 i_1324 (.A1(n_2195), .A2(n_2234), .A3(n_2144), .ZN(n_2194));
   NAND2_X1 i_1325 (.A1(n_1646), .A2(n_1617), .ZN(n_2144));
   NAND2_X1 i_1326 (.A1(n_2197), .A2(n_2196), .ZN(n_2195));
   NOR2_X1 i_1327 (.A1(n_2187), .A2(n_2186), .ZN(n_2196));
   OAI211_X1 i_1328 (.A(n_2224), .B(n_2148), .C1(n_2199), .C2(n_2232), .ZN(
      n_2197));
   AOI21_X1 i_1329 (.A(n_2214), .B1(n_2206), .B2(n_2220), .ZN(n_2199));
   OAI21_X1 i_1330 (.A(n_2209), .B1(n_2052), .B2(n_2479), .ZN(n_2206));
   AOI21_X1 i_1331 (.A(n_2460), .B1(n_2484), .B2(n_2467), .ZN(n_2052));
   INV_X1 i_1332 (.A(n_2453), .ZN(n_2209));
   INV_X1 i_1333 (.A(n_2446), .ZN(n_2214));
   INV_X1 i_1334 (.A(n_2471), .ZN(n_2220));
   NAND2_X1 i_1340 (.A1(n_1584), .A2(n_1551), .ZN(n_2148));
   NAND2_X1 i_1342 (.A1(n_1585), .A2(n_1616), .ZN(n_2224));
   NOR2_X1 i_1343 (.A1(n_1584), .A2(n_1551), .ZN(n_2232));
   INV_X1 i_1346 (.A(n_2080), .ZN(n_2234));
   NAND2_X1 i_1347 (.A1(n_2235), .A2(n_2243), .ZN(out31[52]));
   NAND2_X1 i_1348 (.A1(n_2238), .A2(n_2379), .ZN(n_2235));
   OAI21_X1 i_1350 (.A(n_2245), .B1(n_1725), .B2(n_1746), .ZN(n_2238));
   OAI211_X1 i_1351 (.A(n_2245), .B(n_2378), .C1(n_1725), .C2(n_1746), .ZN(
      n_2243));
   NAND2_X1 i_1352 (.A1(n_2247), .A2(n_2122), .ZN(n_2245));
   INV_X1 i_1354 (.A(n_2253), .ZN(n_2247));
   NAND2_X1 i_1356 (.A1(n_2315), .A2(n_2125), .ZN(n_2253));
   NAND2_X1 i_1357 (.A1(n_2316), .A2(n_2377), .ZN(n_2315));
   OAI21_X1 i_1358 (.A(n_2126), .B1(n_2133), .B2(n_2374), .ZN(n_2316));
   NAND2_X1 i_1359 (.A1(n_1675), .A2(n_1700), .ZN(n_2126));
   NOR2_X1 i_1361 (.A1(n_1675), .A2(n_1700), .ZN(n_2374));
   INV_X1 i_1362 (.A(n_2131), .ZN(n_2377));
   NAND2_X1 i_1364 (.A1(n_1746), .A2(n_1725), .ZN(n_2122));
   INV_X1 i_1366 (.A(n_2379), .ZN(n_2378));
   NOR2_X1 i_1367 (.A1(n_2123), .A2(n_2132), .ZN(n_2379));
   XNOR2_X1 i_1368 (.A(n_2395), .B(n_2384), .ZN(out31[55]));
   NAND2_X1 i_1369 (.A1(n_2381), .A2(n_2387), .ZN(out31[56]));
   OAI21_X1 i_1370 (.A(n_2392), .B1(n_2383), .B2(n_2399), .ZN(n_2381));
   NOR2_X1 i_1372 (.A1(n_2395), .A2(n_2384), .ZN(n_2383));
   NAND2_X1 i_1373 (.A1(n_2084), .A2(n_2107), .ZN(n_2384));
   OAI211_X1 i_1375 (.A(n_2107), .B(n_2391), .C1(n_2395), .C2(n_2400), .ZN(
      n_2387));
   INV_X1 i_1377 (.A(n_2392), .ZN(n_2391));
   AND2_X1 i_1378 (.A1(n_2394), .A2(n_2393), .ZN(n_2392));
   NAND2_X1 i_1379 (.A1(n_1826), .A2(n_1815), .ZN(n_2393));
   INV_X1 i_1380 (.A(n_2112), .ZN(n_2394));
   AOI21_X1 i_1381 (.A(n_2110), .B1(n_2396), .B2(n_2101), .ZN(n_2395));
   AOI21_X1 i_1382 (.A(n_2398), .B1(n_2439), .B2(n_2397), .ZN(n_2396));
   INV_X1 i_1383 (.A(n_2105), .ZN(n_2397));
   INV_X1 i_1384 (.A(n_2102), .ZN(n_2398));
   NAND2_X1 i_1385 (.A1(n_1785), .A2(n_1800), .ZN(n_2101));
   NOR2_X1 i_1386 (.A1(n_1785), .A2(n_1800), .ZN(n_2110));
   INV_X1 i_1387 (.A(n_2399), .ZN(n_2107));
   NOR2_X1 i_1388 (.A1(n_1814), .A2(n_1801), .ZN(n_2399));
   INV_X1 i_1397 (.A(n_2084), .ZN(n_2400));
   XNOR2_X1 i_1449 (.A(n_2419), .B(n_2053), .ZN(out31[58]));
   NAND2_X1 i_1450 (.A1(n_2402), .A2(n_2401), .ZN(out31[59]));
   NAND2_X1 i_1457 (.A1(n_2404), .A2(n_2410), .ZN(n_2401));
   NAND2_X1 i_1459 (.A1(n_2403), .A2(n_2409), .ZN(n_2402));
   INV_X1 i_1461 (.A(n_2404), .ZN(n_2403));
   OAI22_X1 i_1508 (.A1(n_2419), .A2(n_2405), .B1(n_2408), .B2(n_2407), .ZN(
      n_2404));
   INV_X1 i_1510 (.A(n_2406), .ZN(n_2405));
   NAND2_X1 i_1511 (.A1(n_1844), .A2(n_1837), .ZN(n_2406));
   INV_X1 i_1512 (.A(n_2051), .ZN(n_2407));
   INV_X1 i_1513 (.A(n_2049), .ZN(n_2408));
   INV_X1 i_1514 (.A(n_2410), .ZN(n_2409));
   AND2_X1 i_1515 (.A1(n_2411), .A2(n_2090), .ZN(n_2410));
   INV_X1 i_1517 (.A(n_2116), .ZN(n_2411));
   NOR2_X1 i_1518 (.A1(n_2412), .A2(n_2414), .ZN(out31[60]));
   INV_X1 i_1520 (.A(n_2413), .ZN(n_2412));
   NAND3_X1 i_1521 (.A1(n_2417), .A2(n_2090), .A3(n_2415), .ZN(n_2413));
   AOI21_X1 i_1525 (.A(n_2415), .B1(n_2417), .B2(n_2090), .ZN(n_2414));
   INV_X1 i_1526 (.A(n_2416), .ZN(n_2415));
   AOI21_X1 i_1527 (.A(n_2118), .B1(n_1851), .B2(n_1854), .ZN(n_2416));
   NAND2_X1 i_1528 (.A1(n_1850), .A2(n_1845), .ZN(n_2090));
   OAI21_X1 i_1529 (.A(n_2418), .B1(n_2419), .B2(n_2053), .ZN(n_2417));
   NOR2_X1 i_1530 (.A1(n_2117), .A2(n_2116), .ZN(n_2418));
   AOI21_X1 i_1531 (.A(n_2424), .B1(n_2422), .B2(n_2420), .ZN(n_2419));
   INV_X1 i_1532 (.A(n_2421), .ZN(n_2420));
   NAND2_X1 i_1533 (.A1(n_2097), .A2(n_2095), .ZN(n_2421));
   NAND2_X1 i_1534 (.A1(n_2439), .A2(n_2423), .ZN(n_2422));
   INV_X1 i_1535 (.A(n_2085), .ZN(n_2423));
   INV_X1 i_1536 (.A(n_2083), .ZN(n_2424));
   XNOR2_X1 i_1537 (.A(n_2426), .B(n_2425), .ZN(out31[61]));
   NAND2_X1 i_1538 (.A1(n_2089), .A2(n_2086), .ZN(n_2425));
   NAND2_X1 i_1539 (.A1(n_2438), .A2(n_2437), .ZN(n_2426));
   OR2_X1 i_1540 (.A1(n_2428), .A2(n_2427), .ZN(out31[62]));
   AOI21_X1 i_1541 (.A(n_2087), .B1(n_2436), .B2(n_2507), .ZN(n_2427));
   INV_X1 i_1542 (.A(n_2429), .ZN(n_2428));
   NAND3_X1 i_1543 (.A1(n_2436), .A2(n_2087), .A3(n_2507), .ZN(n_2429));
   NAND2_X1 i_1544 (.A1(n_2432), .A2(n_2430), .ZN(out31[63]));
   NAND3_X1 i_1545 (.A1(n_2435), .A2(n_2509), .A3(n_2431), .ZN(n_2430));
   INV_X1 i_1546 (.A(n_2433), .ZN(n_2431));
   NAND2_X1 i_1547 (.A1(n_2434), .A2(n_2433), .ZN(n_2432));
   XOR2_X1 i_1548 (.A(p_30[63]), .B(n_2318), .Z(n_2433));
   NAND2_X1 i_1549 (.A1(n_2435), .A2(n_2509), .ZN(n_2434));
   NAND3_X1 i_1550 (.A1(n_2436), .A2(n_2508), .A3(n_2507), .ZN(n_2435));
   NAND3_X1 i_1551 (.A1(n_2438), .A2(n_2089), .A3(n_2437), .ZN(n_2436));
   AOI21_X1 i_1552 (.A(n_1924), .B1(n_1930), .B2(n_1939), .ZN(n_2437));
   NAND4_X1 i_1553 (.A1(n_2439), .A2(n_1939), .A3(n_1948), .A4(n_2025), .ZN(
      n_2438));
   OAI21_X1 i_1554 (.A(n_2506), .B1(n_2133), .B2(n_2440), .ZN(n_2439));
   NAND2_X1 i_1555 (.A1(n_2029), .A2(n_2441), .ZN(n_2440));
   OR2_X1 i_1556 (.A1(n_1675), .A2(n_1700), .ZN(n_2441));
   AOI21_X1 i_1557 (.A(n_2442), .B1(n_2484), .B2(n_2465), .ZN(n_2133));
   NAND3_X1 i_1558 (.A1(n_2452), .A2(n_2459), .A3(n_2443), .ZN(n_2442));
   INV_X1 i_1559 (.A(n_2444), .ZN(n_2443));
   OAI211_X1 i_1560 (.A(n_2451), .B(n_2445), .C1(n_2446), .C2(n_2477), .ZN(
      n_2444));
   NAND2_X1 i_1561 (.A1(n_1674), .A2(n_1647), .ZN(n_2445));
   AOI21_X1 i_1562 (.A(n_2447), .B1(n_2450), .B2(n_2472), .ZN(n_2446));
   OAI21_X1 i_1563 (.A(n_2449), .B1(n_2448), .B2(n_2473), .ZN(n_2447));
   NAND2_X1 i_1564 (.A1(n_1514), .A2(n_1477), .ZN(n_2448));
   NAND2_X1 i_1565 (.A1(n_1550), .A2(n_1515), .ZN(n_2449));
   NAND2_X1 i_1566 (.A1(n_2140), .A2(n_2139), .ZN(n_2450));
   NAND2_X1 i_1567 (.A1(n_1476), .A2(n_1437), .ZN(n_2139));
   NAND2_X1 i_1568 (.A1(n_1436), .A2(n_1395), .ZN(n_2140));
   INV_X1 i_1569 (.A(n_2142), .ZN(n_2451));
   NAND2_X1 i_1570 (.A1(n_2453), .A2(n_2469), .ZN(n_2452));
   OAI211_X1 i_1571 (.A(n_2455), .B(n_2454), .C1(n_2458), .C2(n_2457), .ZN(
      n_2453));
   OAI211_X1 i_1572 (.A(n_1350), .B(n_1305), .C1(n_1351), .C2(n_1394), .ZN(
      n_2454));
   NAND2_X1 i_1573 (.A1(n_2480), .A2(n_2456), .ZN(n_2455));
   NAND2_X1 i_1574 (.A1(n_2153), .A2(n_2154), .ZN(n_2456));
   NAND2_X1 i_1575 (.A1(n_1256), .A2(n_1207), .ZN(n_2154));
   NAND2_X1 i_1576 (.A1(n_1304), .A2(n_1257), .ZN(n_2153));
   INV_X1 i_1577 (.A(n_1394), .ZN(n_2457));
   INV_X1 i_1578 (.A(n_1351), .ZN(n_2458));
   NAND3_X1 i_1579 (.A1(n_2478), .A2(n_2469), .A3(n_2460), .ZN(n_2459));
   OAI211_X1 i_1580 (.A(n_2462), .B(n_2461), .C1(n_2468), .C2(n_2464), .ZN(
      n_2460));
   NAND2_X1 i_1581 (.A1(n_1206), .A2(n_1155), .ZN(n_2461));
   OR2_X1 i_1582 (.A1(n_2463), .A2(n_2171), .ZN(n_2462));
   NAND2_X1 i_1583 (.A1(n_1154), .A2(n_1101), .ZN(n_2463));
   AND2_X1 i_1584 (.A1(n_2161), .A2(n_2160), .ZN(n_2464));
   NAND2_X1 i_1585 (.A1(n_1100), .A2(n_1045), .ZN(n_2160));
   NAND2_X1 i_1586 (.A1(n_1044), .A2(n_987), .ZN(n_2161));
   INV_X1 i_1587 (.A(n_2466), .ZN(n_2465));
   NAND3_X1 i_1588 (.A1(n_2478), .A2(n_2469), .A3(n_2467), .ZN(n_2466));
   NOR2_X1 i_1589 (.A1(n_2164), .A2(n_2468), .ZN(n_2467));
   OR3_X1 i_1590 (.A1(n_2169), .A2(n_2167), .A3(n_2171), .ZN(n_2468));
   NOR2_X1 i_1591 (.A1(n_1206), .A2(n_1155), .ZN(n_2171));
   NOR2_X1 i_1592 (.A1(n_1100), .A2(n_1045), .ZN(n_2169));
   NOR2_X1 i_1593 (.A1(n_1154), .A2(n_1101), .ZN(n_2167));
   INV_X1 i_1594 (.A(n_2470), .ZN(n_2469));
   OR2_X1 i_1595 (.A1(n_2471), .A2(n_2477), .ZN(n_2470));
   NAND2_X1 i_1596 (.A1(n_2476), .A2(n_2472), .ZN(n_2471));
   NOR3_X1 i_1597 (.A1(n_2474), .A2(n_2475), .A3(n_2473), .ZN(n_2472));
   NOR2_X1 i_1598 (.A1(n_1550), .A2(n_1515), .ZN(n_2473));
   NOR2_X1 i_1599 (.A1(n_1476), .A2(n_1437), .ZN(n_2474));
   NOR2_X1 i_1600 (.A1(n_1514), .A2(n_1477), .ZN(n_2475));
   OR2_X1 i_1601 (.A1(n_1436), .A2(n_1395), .ZN(n_2476));
   OAI21_X1 i_1602 (.A(n_2184), .B1(n_1551), .B2(n_1584), .ZN(n_2477));
   INV_X1 i_1603 (.A(n_2479), .ZN(n_2478));
   OAI21_X1 i_1604 (.A(n_2480), .B1(n_1207), .B2(n_1256), .ZN(n_2479));
   AOI21_X1 i_1605 (.A(n_2481), .B1(n_2483), .B2(n_2482), .ZN(n_2480));
   OAI22_X1 i_1606 (.A1(n_1394), .A2(n_1351), .B1(n_1257), .B2(n_1304), .ZN(
      n_2481));
   INV_X1 i_1607 (.A(n_1350), .ZN(n_2482));
   INV_X1 i_1608 (.A(n_1305), .ZN(n_2483));
   NAND3_X1 i_1609 (.A1(n_2491), .A2(n_2485), .A3(n_2495), .ZN(n_2484));
   NAND4_X1 i_1610 (.A1(n_2252), .A2(n_2504), .A3(n_2490), .A4(n_2486), .ZN(
      n_2485));
   NAND2_X1 i_1611 (.A1(n_2200), .A2(n_2487), .ZN(n_2486));
   NAND2_X1 i_1612 (.A1(n_2488), .A2(n_2489), .ZN(n_2487));
   AOI21_X1 i_1613 (.A(n_2255), .B1(n_2054), .B2(n_2033), .ZN(n_2488));
   INV_X1 i_1614 (.A(n_2262), .ZN(n_2489));
   NOR2_X1 i_1615 (.A1(n_2236), .A2(n_2246), .ZN(n_2490));
   NAND2_X1 i_1616 (.A1(n_2492), .A2(n_2252), .ZN(n_2491));
   NAND2_X1 i_1617 (.A1(n_2493), .A2(n_2208), .ZN(n_2492));
   NAND2_X1 i_1618 (.A1(n_928), .A2(n_869), .ZN(n_2208));
   NAND2_X1 i_1619 (.A1(n_986), .A2(n_2494), .ZN(n_2493));
   INV_X1 i_1620 (.A(n_2328), .ZN(n_2494));
   NAND3_X1 i_1621 (.A1(n_2252), .A2(n_2504), .A3(n_2496), .ZN(n_2495));
   OAI211_X1 i_1622 (.A(n_2503), .B(n_2497), .C1(n_2498), .C2(n_2246), .ZN(
      n_2496));
   NAND2_X1 i_1623 (.A1(n_810), .A2(n_755), .ZN(n_2497));
   INV_X1 i_1624 (.A(n_2499), .ZN(n_2498));
   AOI21_X1 i_1625 (.A(n_2244), .B1(n_2501), .B2(n_2500), .ZN(n_2499));
   AOI22_X1 i_1626 (.A1(n_754), .A2(n_701), .B1(n_649), .B2(n_700), .ZN(n_2500));
   NAND3_X1 i_1627 (.A1(n_2502), .A2(n_2239), .A3(n_2241), .ZN(n_2501));
   NAND2_X1 i_1628 (.A1(n_2217), .A2(n_2216), .ZN(n_2502));
   INV_X1 i_1629 (.A(n_2242), .ZN(n_2241));
   INV_X1 i_1630 (.A(n_2240), .ZN(n_2239));
   NOR2_X1 i_1631 (.A1(n_754), .A2(n_701), .ZN(n_2244));
   NOR2_X1 i_1632 (.A1(n_810), .A2(n_755), .ZN(n_2246));
   INV_X1 i_1633 (.A(n_2210), .ZN(n_2503));
   NOR2_X1 i_1634 (.A1(n_2249), .A2(n_2251), .ZN(n_2504));
   NOR2_X1 i_1635 (.A1(n_868), .A2(n_811), .ZN(n_2251));
   NOR2_X1 i_1636 (.A1(n_928), .A2(n_869), .ZN(n_2249));
   NAND2_X1 i_1637 (.A1(n_2327), .A2(n_2505), .ZN(n_2252));
   INV_X1 i_1638 (.A(n_986), .ZN(n_2327));
   INV_X1 i_1639 (.A(n_929), .ZN(n_2505));
   INV_X1 i_1640 (.A(n_2088), .ZN(n_2506));
   OR2_X1 i_1641 (.A1(n_1856), .A2(n_1855), .ZN(n_2507));
   OR2_X1 i_1642 (.A1(n_1857), .A2(n_2043), .ZN(n_2508));
   NAND2_X1 i_1643 (.A1(n_1857), .A2(n_2043), .ZN(n_2509));
endmodule

module datapath__0_65(p_0, in2);
   output [31:0]p_0;
   input [31:0]in2;

   AOI21_X1 i_0 (.A(n_62), .B1(in2[1]), .B2(in2[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_60), .B1(in2[2]), .B2(n_61), .ZN(p_0[2]));
   AOI21_X1 i_3 (.A(n_5), .B1(in2[4]), .B2(n_57), .ZN(p_0[4]));
   XNOR2_X1 i_67 (.A(in2[31]), .B(n_37), .ZN(p_0[31]));
   INV_X1 i_2 (.A(n_59), .ZN(n_60));
   NOR2_X1 i_4 (.A1(in2[28]), .A2(in2[29]), .ZN(n_0));
   NAND4_X1 i_5 (.A1(n_100), .A2(n_104), .A3(n_101), .A4(n_0), .ZN(n_1));
   INV_X1 i_6 (.A(n_1), .ZN(n_2));
   INV_X1 i_7 (.A(n_105), .ZN(n_3));
   AOI21_X1 i_8 (.A(n_2), .B1(n_3), .B2(in2[29]), .ZN(p_0[29]));
   NAND4_X1 i_9 (.A1(n_100), .A2(n_104), .A3(n_0), .A4(n_101), .ZN(n_4));
   NOR2_X1 i_10 (.A1(n_4), .A2(in2[30]), .ZN(n_6));
   AOI21_X1 i_11 (.A(n_6), .B1(n_1), .B2(in2[30]), .ZN(p_0[30]));
   BUF_X1 i_12 (.A(n_96), .Z(n_57));
   BUF_X1 i_13 (.A(n_97), .Z(n_5));
   BUF_X1 i_14 (.A(n_6), .Z(n_37));
   INV_X1 i_15 (.A(in2[20]), .ZN(n_7));
   OR3_X1 i_16 (.A1(n_102), .A2(n_98), .A3(n_99), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_103), .B1(n_8), .B2(in2[21]), .ZN(p_0[21]));
   NOR4_X1 i_18 (.A1(in2[3]), .A2(in2[0]), .A3(in2[2]), .A4(in2[1]), .ZN(n_9));
   INV_X1 i_19 (.A(n_9), .ZN(n_10));
   NOR2_X1 i_20 (.A1(in2[0]), .A2(in2[1]), .ZN(n_11));
   INV_X1 i_21 (.A(n_11), .ZN(n_12));
   OR2_X1 i_22 (.A1(n_12), .A2(in2[2]), .ZN(n_13));
   AOI21_X1 i_23 (.A(n_9), .B1(n_13), .B2(in2[3]), .ZN(p_0[3]));
   NOR2_X1 i_24 (.A1(n_10), .A2(in2[4]), .ZN(n_14));
   INV_X1 i_25 (.A(n_14), .ZN(n_15));
   NOR2_X1 i_26 (.A1(n_15), .A2(in2[5]), .ZN(n_16));
   AOI21_X1 i_27 (.A(n_16), .B1(n_15), .B2(in2[5]), .ZN(p_0[5]));
   NOR3_X1 i_28 (.A1(n_15), .A2(in2[5]), .A3(in2[6]), .ZN(n_17));
   INV_X1 i_29 (.A(n_16), .ZN(n_18));
   AOI21_X1 i_30 (.A(n_17), .B1(n_18), .B2(in2[6]), .ZN(p_0[6]));
   NOR4_X1 i_31 (.A1(in2[4]), .A2(in2[5]), .A3(in2[6]), .A4(in2[7]), .ZN(n_19));
   INV_X1 i_32 (.A(n_19), .ZN(n_20));
   NOR2_X1 i_33 (.A1(n_10), .A2(n_20), .ZN(n_21));
   INV_X1 i_34 (.A(n_21), .ZN(n_22));
   INV_X1 i_35 (.A(n_17), .ZN(n_23));
   AOI21_X1 i_36 (.A(n_21), .B1(n_23), .B2(in2[7]), .ZN(p_0[7]));
   XNOR2_X1 i_37 (.A(n_21), .B(in2[8]), .ZN(p_0[8]));
   NOR3_X1 i_38 (.A1(n_22), .A2(in2[8]), .A3(in2[9]), .ZN(n_24));
   OR2_X1 i_39 (.A1(n_22), .A2(in2[8]), .ZN(n_25));
   AOI21_X1 i_40 (.A(n_24), .B1(n_25), .B2(in2[9]), .ZN(p_0[9]));
   NOR4_X1 i_41 (.A1(n_10), .A2(n_20), .A3(in2[10]), .A4(in2[8]), .ZN(n_26));
   INV_X1 i_42 (.A(in2[9]), .ZN(n_27));
   NAND2_X1 i_43 (.A1(n_26), .A2(n_27), .ZN(n_28));
   INV_X1 i_44 (.A(n_28), .ZN(n_29));
   INV_X1 i_45 (.A(n_24), .ZN(n_30));
   AOI21_X1 i_46 (.A(n_29), .B1(n_30), .B2(in2[10]), .ZN(p_0[10]));
   NOR4_X1 i_47 (.A1(in2[8]), .A2(in2[9]), .A3(in2[10]), .A4(in2[11]), .ZN(n_31));
   INV_X1 i_48 (.A(n_31), .ZN(n_32));
   NOR3_X1 i_49 (.A1(n_10), .A2(n_20), .A3(n_32), .ZN(n_33));
   AOI21_X1 i_50 (.A(n_33), .B1(n_28), .B2(in2[11]), .ZN(p_0[11]));
   NOR4_X1 i_51 (.A1(n_32), .A2(n_10), .A3(n_20), .A4(in2[12]), .ZN(n_34));
   INV_X1 i_52 (.A(n_33), .ZN(n_35));
   AOI21_X1 i_53 (.A(n_34), .B1(n_35), .B2(in2[12]), .ZN(p_0[12]));
   INV_X1 i_54 (.A(n_34), .ZN(n_36));
   NOR2_X1 i_55 (.A1(n_36), .A2(in2[13]), .ZN(n_38));
   AOI21_X1 i_56 (.A(n_38), .B1(n_36), .B2(in2[13]), .ZN(p_0[13]));
   NOR4_X1 i_57 (.A1(n_35), .A2(in2[12]), .A3(in2[13]), .A4(in2[14]), .ZN(n_39));
   INV_X1 i_58 (.A(n_38), .ZN(n_40));
   AOI21_X1 i_59 (.A(n_39), .B1(n_40), .B2(in2[14]), .ZN(p_0[14]));
   NOR4_X1 i_60 (.A1(in2[12]), .A2(in2[13]), .A3(in2[14]), .A4(in2[15]), 
      .ZN(n_41));
   NAND4_X1 i_61 (.A1(n_9), .A2(n_19), .A3(n_31), .A4(n_41), .ZN(n_42));
   INV_X1 i_62 (.A(n_42), .ZN(n_43));
   INV_X1 i_63 (.A(n_39), .ZN(n_44));
   AOI21_X1 i_64 (.A(n_43), .B1(n_44), .B2(in2[15]), .ZN(p_0[15]));
   INV_X1 i_65 (.A(n_41), .ZN(n_45));
   NOR4_X1 i_66 (.A1(n_22), .A2(in2[16]), .A3(n_32), .A4(n_45), .ZN(n_46));
   AOI21_X1 i_68 (.A(n_46), .B1(n_42), .B2(in2[16]), .ZN(p_0[16]));
   NOR4_X1 i_69 (.A1(n_35), .A2(in2[16]), .A3(in2[17]), .A4(n_45), .ZN(n_47));
   INV_X1 i_70 (.A(n_46), .ZN(n_48));
   AOI21_X1 i_71 (.A(n_47), .B1(n_48), .B2(in2[17]), .ZN(p_0[17]));
   NOR4_X1 i_72 (.A1(n_35), .A2(in2[18]), .A3(in2[17]), .A4(n_45), .ZN(n_49));
   INV_X1 i_73 (.A(in2[16]), .ZN(n_50));
   NAND2_X1 i_74 (.A1(n_49), .A2(n_50), .ZN(n_51));
   INV_X1 i_75 (.A(n_51), .ZN(n_52));
   INV_X1 i_76 (.A(n_47), .ZN(n_53));
   AOI21_X1 i_77 (.A(n_52), .B1(n_53), .B2(in2[18]), .ZN(p_0[18]));
   NOR4_X1 i_78 (.A1(n_32), .A2(in2[17]), .A3(in2[18]), .A4(in2[19]), .ZN(n_54));
   NAND2_X1 i_79 (.A1(n_54), .A2(n_50), .ZN(n_55));
   NOR3_X1 i_80 (.A1(n_10), .A2(n_20), .A3(n_45), .ZN(n_56));
   INV_X1 i_81 (.A(n_56), .ZN(n_58));
   NOR2_X1 i_82 (.A1(n_55), .A2(n_58), .ZN(n_63));
   AOI21_X1 i_83 (.A(n_63), .B1(n_51), .B2(in2[19]), .ZN(p_0[19]));
   NOR3_X1 i_84 (.A1(n_55), .A2(n_58), .A3(in2[20]), .ZN(n_64));
   INV_X1 i_85 (.A(n_63), .ZN(n_65));
   AOI21_X1 i_86 (.A(n_64), .B1(n_65), .B2(in2[20]), .ZN(p_0[20]));
   NOR3_X1 i_87 (.A1(in2[20]), .A2(in2[22]), .A3(in2[21]), .ZN(n_66));
   NAND2_X1 i_88 (.A1(n_41), .A2(n_7), .ZN(n_67));
   OR4_X1 i_89 (.A1(n_55), .A2(n_10), .A3(n_20), .A4(n_67), .ZN(n_68));
   NOR2_X1 i_90 (.A1(n_68), .A2(in2[21]), .ZN(n_69));
   INV_X1 i_91 (.A(n_66), .ZN(n_70));
   OR2_X1 i_92 (.A1(in2[18]), .A2(in2[19]), .ZN(n_71));
   OR2_X1 i_93 (.A1(in2[16]), .A2(in2[17]), .ZN(n_72));
   NOR3_X1 i_94 (.A1(n_70), .A2(n_71), .A3(n_72), .ZN(n_73));
   NAND4_X1 i_95 (.A1(n_21), .A2(n_31), .A3(n_41), .A4(n_73), .ZN(n_74));
   INV_X1 i_96 (.A(n_74), .ZN(n_75));
   INV_X1 i_97 (.A(n_69), .ZN(n_76));
   AOI21_X1 i_98 (.A(n_75), .B1(n_76), .B2(in2[22]), .ZN(p_0[22]));
   NOR4_X1 i_99 (.A1(n_70), .A2(n_72), .A3(n_71), .A4(in2[23]), .ZN(n_77));
   INV_X1 i_100 (.A(n_77), .ZN(n_78));
   NOR2_X1 i_101 (.A1(n_42), .A2(n_78), .ZN(n_79));
   AOI21_X1 i_102 (.A(n_79), .B1(n_74), .B2(in2[23]), .ZN(p_0[23]));
   NOR4_X1 i_103 (.A1(n_35), .A2(n_78), .A3(in2[24]), .A4(n_45), .ZN(n_80));
   INV_X1 i_104 (.A(n_79), .ZN(n_81));
   AOI21_X1 i_105 (.A(n_80), .B1(n_81), .B2(in2[24]), .ZN(p_0[24]));
   NOR3_X1 i_106 (.A1(in2[23]), .A2(in2[24]), .A3(in2[25]), .ZN(n_82));
   AND4_X1 i_107 (.A1(n_33), .A2(n_73), .A3(n_41), .A4(n_82), .ZN(n_83));
   INV_X1 i_108 (.A(n_80), .ZN(n_84));
   AOI21_X1 i_109 (.A(n_83), .B1(n_84), .B2(in2[25]), .ZN(p_0[25]));
   NOR3_X1 i_110 (.A1(in2[24]), .A2(in2[25]), .A3(in2[26]), .ZN(n_85));
   NAND4_X1 i_111 (.A1(n_77), .A2(n_33), .A3(n_41), .A4(n_85), .ZN(n_86));
   INV_X1 i_112 (.A(n_86), .ZN(n_87));
   INV_X1 i_113 (.A(n_55), .ZN(n_88));
   NAND4_X1 i_114 (.A1(n_88), .A2(n_66), .A3(n_56), .A4(n_82), .ZN(n_89));
   AOI21_X1 i_115 (.A(n_87), .B1(n_89), .B2(in2[26]), .ZN(p_0[26]));
   NOR2_X1 i_116 (.A1(in2[23]), .A2(in2[27]), .ZN(n_90));
   AND2_X1 i_117 (.A1(n_85), .A2(n_90), .ZN(n_91));
   NAND4_X1 i_118 (.A1(n_33), .A2(n_41), .A3(n_73), .A4(n_91), .ZN(n_92));
   INV_X1 i_119 (.A(n_92), .ZN(n_93));
   AOI21_X1 i_120 (.A(n_93), .B1(n_86), .B2(in2[27]), .ZN(p_0[27]));
   NAND4_X1 i_121 (.A1(n_88), .A2(n_85), .A3(n_56), .A4(n_90), .ZN(n_94));
   NOR3_X1 i_122 (.A1(n_94), .A2(in2[28]), .A3(n_70), .ZN(n_95));
   AOI21_X1 i_123 (.A(n_95), .B1(n_92), .B2(in2[28]), .ZN(p_0[28]));
   BUF_X1 i_124 (.A(n_10), .Z(n_96));
   BUF_X1 i_125 (.A(n_12), .Z(n_61));
   BUF_X1 i_126 (.A(n_11), .Z(n_62));
   BUF_X1 i_127 (.A(n_13), .Z(n_59));
   BUF_X1 i_128 (.A(n_14), .Z(n_97));
   BUF_X1 i_129 (.A(n_22), .Z(n_98));
   BUF_X1 i_130 (.A(n_55), .Z(n_99));
   BUF_X1 i_131 (.A(n_63), .Z(n_100));
   BUF_X1 i_132 (.A(n_66), .Z(n_101));
   BUF_X1 i_133 (.A(n_67), .Z(n_102));
   BUF_X1 i_134 (.A(n_69), .Z(n_103));
   BUF_X1 i_135 (.A(n_91), .Z(n_104));
   BUF_X1 i_136 (.A(n_95), .Z(n_105));
endmodule

module datapath(p_0, in1);
   output [31:0]p_0;
   input [31:0]in1;

   AOI21_X1 i_0 (.A(n_80), .B1(in1[1]), .B2(in1[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_7), .B1(in1[2]), .B2(n_79), .ZN(p_0[2]));
   AOI21_X1 i_2 (.A(n_82), .B1(in1[4]), .B2(n_77), .ZN(p_0[4]));
   AOI21_X1 i_3 (.A(n_6), .B1(in1[7]), .B2(n_0), .ZN(p_0[7]));
   INV_X1 i_4 (.A(n_78), .ZN(n_0));
   AOI21_X1 i_5 (.A(n_2), .B1(in1[30]), .B2(n_1), .ZN(p_0[30]));
   INV_X1 i_6 (.A(n_3), .ZN(n_1));
   XNOR2_X1 i_7 (.A(in1[31]), .B(n_2), .ZN(p_0[31]));
   NOR4_X1 i_8 (.A1(in1[29]), .A2(in1[28]), .A3(in1[30]), .A4(n_4), .ZN(n_2));
   INV_X1 i_9 (.A(n_87), .ZN(n_3));
   NAND2_X1 i_10 (.A1(n_84), .A2(n_86), .ZN(n_4));
   NAND3_X1 i_11 (.A1(n_27), .A2(n_24), .A3(n_22), .ZN(n_5));
   INV_X1 i_12 (.A(n_83), .ZN(n_6));
   INV_X1 i_13 (.A(n_81), .ZN(n_7));
   INV_X1 i_14 (.A(in1[29]), .ZN(n_8));
   OR2_X1 i_15 (.A1(n_10), .A2(in1[27]), .ZN(n_9));
   NAND3_X1 i_16 (.A1(n_11), .A2(n_62), .A3(n_85), .ZN(n_10));
   INV_X1 i_17 (.A(in1[26]), .ZN(n_11));
   NAND3_X1 i_18 (.A1(n_15), .A2(n_14), .A3(n_13), .ZN(n_12));
   INV_X1 i_19 (.A(in1[20]), .ZN(n_13));
   INV_X1 i_20 (.A(in1[21]), .ZN(n_14));
   INV_X1 i_21 (.A(in1[22]), .ZN(n_15));
   NOR4_X1 i_22 (.A1(in1[2]), .A2(in1[0]), .A3(in1[1]), .A4(in1[3]), .ZN(n_16));
   INV_X1 i_23 (.A(n_16), .ZN(n_17));
   NOR2_X1 i_24 (.A1(n_17), .A2(n_5), .ZN(n_18));
   NOR2_X1 i_25 (.A1(in1[0]), .A2(in1[1]), .ZN(n_19));
   INV_X1 i_26 (.A(n_19), .ZN(n_20));
   OR2_X1 i_27 (.A1(n_20), .A2(in1[2]), .ZN(n_21));
   AOI21_X1 i_28 (.A(n_16), .B1(n_21), .B2(in1[3]), .ZN(p_0[3]));
   INV_X1 i_29 (.A(in1[4]), .ZN(n_22));
   NOR2_X1 i_30 (.A1(n_17), .A2(in1[4]), .ZN(n_23));
   INV_X1 i_31 (.A(in1[5]), .ZN(n_24));
   INV_X1 i_32 (.A(n_23), .ZN(n_25));
   NOR2_X1 i_33 (.A1(n_25), .A2(in1[5]), .ZN(n_26));
   AOI21_X1 i_34 (.A(n_26), .B1(n_25), .B2(in1[5]), .ZN(p_0[5]));
   INV_X1 i_35 (.A(in1[6]), .ZN(n_27));
   INV_X1 i_36 (.A(n_26), .ZN(n_28));
   AOI21_X1 i_37 (.A(n_18), .B1(n_28), .B2(in1[6]), .ZN(p_0[6]));
   NOR4_X1 i_38 (.A1(in1[4]), .A2(in1[5]), .A3(in1[6]), .A4(in1[7]), .ZN(n_29));
   NAND2_X1 i_39 (.A1(n_16), .A2(n_29), .ZN(n_30));
   NOR2_X1 i_40 (.A1(n_30), .A2(in1[8]), .ZN(n_31));
   AOI21_X1 i_41 (.A(n_31), .B1(n_30), .B2(in1[8]), .ZN(p_0[8]));
   XNOR2_X1 i_42 (.A(n_31), .B(in1[9]), .ZN(p_0[9]));
   INV_X1 i_43 (.A(n_31), .ZN(n_32));
   NOR3_X1 i_44 (.A1(n_32), .A2(in1[10]), .A3(in1[9]), .ZN(n_33));
   OR2_X1 i_45 (.A1(n_32), .A2(in1[9]), .ZN(n_34));
   AOI21_X1 i_46 (.A(n_33), .B1(n_34), .B2(in1[10]), .ZN(p_0[10]));
   NOR4_X1 i_47 (.A1(in1[8]), .A2(in1[10]), .A3(in1[9]), .A4(in1[11]), .ZN(n_35));
   NAND3_X1 i_48 (.A1(n_16), .A2(n_29), .A3(n_35), .ZN(n_36));
   INV_X1 i_49 (.A(n_36), .ZN(n_37));
   INV_X1 i_50 (.A(n_33), .ZN(n_38));
   AOI21_X1 i_51 (.A(n_37), .B1(n_38), .B2(in1[11]), .ZN(p_0[11]));
   NOR2_X1 i_52 (.A1(n_36), .A2(in1[12]), .ZN(n_39));
   AOI21_X1 i_53 (.A(n_39), .B1(n_36), .B2(in1[12]), .ZN(p_0[12]));
   XNOR2_X1 i_54 (.A(n_39), .B(in1[13]), .ZN(p_0[13]));
   INV_X1 i_55 (.A(n_39), .ZN(n_40));
   NOR3_X1 i_56 (.A1(n_40), .A2(in1[14]), .A3(in1[13]), .ZN(n_41));
   OR2_X1 i_57 (.A1(n_40), .A2(in1[13]), .ZN(n_42));
   AOI21_X1 i_58 (.A(n_41), .B1(n_42), .B2(in1[14]), .ZN(p_0[14]));
   NOR4_X1 i_59 (.A1(in1[12]), .A2(in1[14]), .A3(in1[13]), .A4(in1[15]), 
      .ZN(n_43));
   NAND4_X1 i_60 (.A1(n_16), .A2(n_29), .A3(n_35), .A4(n_43), .ZN(n_44));
   INV_X1 i_61 (.A(n_44), .ZN(n_45));
   INV_X1 i_62 (.A(n_41), .ZN(n_46));
   AOI21_X1 i_63 (.A(n_45), .B1(n_46), .B2(in1[15]), .ZN(p_0[15]));
   NOR2_X1 i_64 (.A1(n_44), .A2(in1[16]), .ZN(n_47));
   AOI21_X1 i_65 (.A(n_47), .B1(n_44), .B2(in1[16]), .ZN(p_0[16]));
   XNOR2_X1 i_66 (.A(n_47), .B(in1[17]), .ZN(p_0[17]));
   NOR4_X1 i_67 (.A1(n_44), .A2(in1[16]), .A3(in1[17]), .A4(in1[18]), .ZN(n_48));
   INV_X1 i_68 (.A(in1[17]), .ZN(n_49));
   NAND2_X1 i_69 (.A1(n_47), .A2(n_49), .ZN(n_50));
   AOI21_X1 i_70 (.A(n_48), .B1(n_50), .B2(in1[18]), .ZN(p_0[18]));
   INV_X1 i_71 (.A(n_43), .ZN(n_51));
   OR4_X1 i_72 (.A1(in1[16]), .A2(in1[17]), .A3(in1[18]), .A4(in1[19]), .ZN(n_52));
   NOR3_X1 i_73 (.A1(n_36), .A2(n_51), .A3(n_52), .ZN(n_53));
   INV_X1 i_74 (.A(n_48), .ZN(n_54));
   AOI21_X1 i_75 (.A(n_53), .B1(n_54), .B2(in1[19]), .ZN(p_0[19]));
   XNOR2_X1 i_76 (.A(n_53), .B(in1[20]), .ZN(p_0[20]));
   INV_X1 i_77 (.A(n_53), .ZN(n_55));
   NOR3_X1 i_78 (.A1(n_55), .A2(in1[20]), .A3(in1[21]), .ZN(n_56));
   OR2_X1 i_79 (.A1(n_55), .A2(in1[20]), .ZN(n_57));
   AOI21_X1 i_80 (.A(n_56), .B1(n_57), .B2(in1[21]), .ZN(p_0[21]));
   NOR4_X1 i_81 (.A1(n_36), .A2(n_12), .A3(n_51), .A4(n_52), .ZN(n_58));
   INV_X1 i_82 (.A(n_56), .ZN(n_59));
   AOI21_X1 i_83 (.A(n_58), .B1(n_59), .B2(in1[22]), .ZN(p_0[22]));
   NOR4_X1 i_84 (.A1(n_44), .A2(n_12), .A3(in1[23]), .A4(n_52), .ZN(n_60));
   INV_X1 i_85 (.A(n_58), .ZN(n_61));
   AOI21_X1 i_86 (.A(n_60), .B1(n_61), .B2(in1[23]), .ZN(p_0[23]));
   XNOR2_X1 i_87 (.A(n_60), .B(in1[24]), .ZN(p_0[24]));
   INV_X1 i_88 (.A(in1[25]), .ZN(n_62));
   INV_X1 i_89 (.A(in1[24]), .ZN(n_63));
   NOR4_X1 i_90 (.A1(n_61), .A2(in1[23]), .A3(in1[25]), .A4(in1[24]), .ZN(n_64));
   NAND2_X1 i_91 (.A1(n_60), .A2(n_63), .ZN(n_65));
   AOI21_X1 i_92 (.A(n_64), .B1(n_65), .B2(in1[25]), .ZN(p_0[25]));
   NOR4_X1 i_93 (.A1(n_55), .A2(n_12), .A3(in1[23]), .A4(n_10), .ZN(n_66));
   INV_X1 i_94 (.A(n_64), .ZN(n_67));
   AOI21_X1 i_95 (.A(n_66), .B1(n_67), .B2(in1[26]), .ZN(p_0[26]));
   INV_X1 i_96 (.A(n_9), .ZN(n_68));
   AND2_X1 i_97 (.A1(n_68), .A2(n_60), .ZN(n_69));
   INV_X1 i_98 (.A(n_66), .ZN(n_70));
   AOI21_X1 i_99 (.A(n_69), .B1(n_70), .B2(in1[27]), .ZN(p_0[27]));
   NOR4_X1 i_100 (.A1(n_61), .A2(in1[23]), .A3(n_9), .A4(in1[28]), .ZN(n_71));
   INV_X1 i_101 (.A(n_69), .ZN(n_72));
   AOI21_X1 i_102 (.A(n_71), .B1(n_72), .B2(in1[28]), .ZN(p_0[28]));
   INV_X1 i_103 (.A(in1[28]), .ZN(n_73));
   NAND4_X1 i_104 (.A1(n_60), .A2(n_68), .A3(n_73), .A4(n_8), .ZN(n_74));
   INV_X1 i_105 (.A(n_74), .ZN(n_75));
   INV_X1 i_106 (.A(n_71), .ZN(n_76));
   AOI21_X1 i_107 (.A(n_75), .B1(n_76), .B2(in1[29]), .ZN(p_0[29]));
   BUF_X1 i_108 (.A(n_17), .Z(n_77));
   BUF_X1 i_109 (.A(n_18), .Z(n_78));
   BUF_X1 i_110 (.A(n_20), .Z(n_79));
   BUF_X1 i_111 (.A(n_19), .Z(n_80));
   BUF_X1 i_112 (.A(n_21), .Z(n_81));
   BUF_X1 i_113 (.A(n_23), .Z(n_82));
   BUF_X1 i_114 (.A(n_30), .Z(n_83));
   BUF_X1 i_115 (.A(n_60), .Z(n_84));
   BUF_X1 i_116 (.A(n_63), .Z(n_85));
   BUF_X1 i_117 (.A(n_68), .Z(n_86));
   BUF_X1 i_118 (.A(n_74), .Z(n_87));
endmodule

module sequential_multiplier(clk, rst, in1, in2, out);
   input clk;
   input rst;
   input [31:0]in1;
   input [31:0]in2;
   output [63:0]out;

   wire n_8_0;
   wire n_8_1;
   wire n_8_2;
   wire n_8_3;
   wire n_8_0_6;
   wire n_8_4;
   wire n_8_5;
   wire n_8_0_8;
   wire n_8_6;
   wire n_8_7;
   wire n_8_0_10;
   wire n_8_8;
   wire n_8_9;
   wire n_8_10;
   wire n_8_11;
   wire n_8_0_14;
   wire n_8_12;
   wire n_8_0_15;
   wire n_8_13;
   wire n_8_0_16;
   wire n_8_14;
   wire n_8_0_17;
   wire n_8_15;
   wire n_8_0_18;
   wire n_8_16;
   wire n_8_0_19;
   wire n_8_17;
   wire n_8_0_20;
   wire n_8_18;
   wire n_8_0_21;
   wire n_8_19;
   wire n_8_0_22;
   wire n_8_20;
   wire n_8_0_23;
   wire n_8_21;
   wire n_8_0_24;
   wire n_8_22;
   wire n_8_23;
   wire n_8_24;
   wire n_8_26;
   wire n_8_29;
   wire n_8_30;
   wire n_8_31;
   wire n_8_0_34;
   wire n_8_32;
   wire n_8_33;
   wire n_8_34;
   wire n_8_35;
   wire n_8_36;
   wire n_8_37;
   wire n_8_38;
   wire n_8_39;
   wire n_8_40;
   wire n_8_41;
   wire n_8_42;
   wire n_8_43;
   wire n_8_44;
   wire n_8_45;
   wire n_8_46;
   wire n_8_47;
   wire n_8_48;
   wire n_8_49;
   wire n_8_50;
   wire n_8_51;
   wire n_8_52;
   wire n_8_53;
   wire n_8_54;
   wire n_8_55;
   wire n_8_56;
   wire n_8_57;
   wire n_8_58;
   wire n_8_59;
   wire n_8_60;
   wire n_8_61;
   wire n_8_62;
   wire n_8_63;
   wire n_8_64;
   wire n_8_66;
   wire n_8_67;
   wire n_8_68;
   wire n_8_69;
   wire n_8_70;
   wire n_8_71;
   wire n_8_72;
   wire n_8_73;
   wire n_8_74;
   wire n_8_75;
   wire n_8_76;
   wire n_8_77;
   wire n_8_78;
   wire n_8_79;
   wire n_8_80;
   wire n_8_81;
   wire n_8_82;
   wire n_8_83;
   wire n_8_84;
   wire n_8_85;
   wire n_8_86;
   wire n_8_87;
   wire n_8_88;
   wire n_8_89;
   wire n_8_90;
   wire n_8_91;
   wire n_8_92;
   wire n_8_93;
   wire n_8_94;
   wire n_8_95;
   wire n_8_96;
   wire n_8_97;
   wire n_8_101;
   wire n_8_102;
   wire n_8_103;
   wire n_8_104;
   wire n_8_105;
   wire n_8_106;
   wire n_8_107;
   wire n_8_108;
   wire n_8_109;
   wire n_8_110;
   wire n_8_111;
   wire n_8_112;
   wire n_8_113;
   wire n_8_114;
   wire n_8_115;
   wire n_8_116;
   wire n_8_117;
   wire n_8_118;
   wire n_8_119;
   wire n_8_120;
   wire n_8_121;
   wire n_8_122;
   wire n_8_123;
   wire n_8_124;
   wire n_8_125;
   wire n_8_126;
   wire n_8_127;
   wire n_8_128;
   wire n_8_129;
   wire n_8_130;
   wire n_8_132;
   wire n_8_134;
   wire n_8_135;
   wire n_8_136;
   wire n_8_137;
   wire n_8_138;
   wire n_8_139;
   wire n_8_140;
   wire n_8_141;
   wire n_8_142;
   wire n_8_143;
   wire n_8_144;
   wire n_8_145;
   wire n_8_146;
   wire n_8_147;
   wire n_8_148;
   wire n_8_149;
   wire n_8_150;
   wire n_8_151;
   wire n_8_152;
   wire n_8_153;
   wire n_8_154;
   wire n_8_155;
   wire n_8_156;
   wire n_8_157;
   wire n_8_158;
   wire n_8_159;
   wire n_8_160;
   wire n_8_161;
   wire n_8_162;
   wire n_8_163;
   wire n_8_165;
   wire n_8_166;
   wire n_8_167;
   wire n_8_168;
   wire n_8_169;
   wire n_8_170;
   wire n_8_171;
   wire n_8_172;
   wire n_8_173;
   wire n_8_174;
   wire n_8_175;
   wire n_8_176;
   wire n_8_177;
   wire n_8_178;
   wire n_8_179;
   wire n_8_180;
   wire n_8_181;
   wire n_8_182;
   wire n_8_183;
   wire n_8_184;
   wire n_8_185;
   wire n_8_186;
   wire n_8_187;
   wire n_8_188;
   wire n_8_189;
   wire n_8_190;
   wire n_8_191;
   wire n_8_192;
   wire n_8_193;
   wire n_8_194;
   wire n_8_195;
   wire n_8_196;
   wire n_8_200;
   wire n_8_201;
   wire n_8_202;
   wire n_8_203;
   wire n_8_204;
   wire n_8_205;
   wire n_8_206;
   wire n_8_207;
   wire n_8_208;
   wire n_8_209;
   wire n_8_210;
   wire n_8_211;
   wire n_8_212;
   wire n_8_213;
   wire n_8_214;
   wire n_8_215;
   wire n_8_216;
   wire n_8_217;
   wire n_8_218;
   wire n_8_219;
   wire n_8_220;
   wire n_8_221;
   wire n_8_222;
   wire n_8_223;
   wire n_8_224;
   wire n_8_225;
   wire n_8_226;
   wire n_8_227;
   wire n_8_228;
   wire n_8_229;
   wire n_8_230;
   wire n_8_235;
   wire n_8_237;
   wire n_8_239;
   wire n_8_243;
   wire n_8_244;
   wire n_8_245;
   wire n_8_246;
   wire n_8_247;
   wire n_8_248;
   wire n_8_249;
   wire n_8_250;
   wire n_8_251;
   wire n_8_252;
   wire n_8_253;
   wire n_8_254;
   wire n_8_255;
   wire n_8_256;
   wire n_8_257;
   wire n_8_258;
   wire n_8_259;
   wire n_8_260;
   wire n_8_261;
   wire n_8_262;
   wire n_8_0_41;
   wire n_8_263;
   wire n_8_264;
   wire n_8_265;
   wire n_8_266;
   wire n_8_267;
   wire n_8_268;
   wire n_8_269;
   wire n_8_270;
   wire n_8_271;
   wire n_8_272;
   wire n_8_273;
   wire n_8_274;
   wire n_8_275;
   wire n_8_276;
   wire n_8_277;
   wire n_8_278;
   wire n_8_279;
   wire n_8_280;
   wire n_8_281;
   wire n_8_282;
   wire n_8_283;
   wire n_8_284;
   wire n_8_285;
   wire n_8_286;
   wire n_8_287;
   wire n_8_288;
   wire n_8_289;
   wire n_8_290;
   wire n_8_291;
   wire n_8_292;
   wire n_8_293;
   wire n_8_294;
   wire n_8_295;
   wire n_8_0_42;
   wire n_8_296;
   wire n_8_297;
   wire n_8_298;
   wire n_8_299;
   wire n_8_300;
   wire n_8_301;
   wire n_8_302;
   wire n_8_303;
   wire n_8_304;
   wire n_8_305;
   wire n_8_306;
   wire n_8_307;
   wire n_8_308;
   wire n_8_309;
   wire n_8_310;
   wire n_8_311;
   wire n_8_312;
   wire n_8_313;
   wire n_8_314;
   wire n_8_315;
   wire n_8_316;
   wire n_8_317;
   wire n_8_318;
   wire n_8_319;
   wire n_8_320;
   wire n_8_321;
   wire n_8_322;
   wire n_8_323;
   wire n_8_324;
   wire n_8_325;
   wire n_8_326;
   wire n_8_327;
   wire n_8_328;
   wire n_8_0_43;
   wire n_8_329;
   wire n_8_330;
   wire n_8_331;
   wire n_8_332;
   wire n_8_333;
   wire n_8_334;
   wire n_8_335;
   wire n_8_336;
   wire n_8_337;
   wire n_8_338;
   wire n_8_339;
   wire n_8_340;
   wire n_8_341;
   wire n_8_342;
   wire n_8_343;
   wire n_8_344;
   wire n_8_345;
   wire n_8_346;
   wire n_8_347;
   wire n_8_348;
   wire n_8_349;
   wire n_8_350;
   wire n_8_351;
   wire n_8_352;
   wire n_8_353;
   wire n_8_354;
   wire n_8_355;
   wire n_8_356;
   wire n_8_357;
   wire n_8_358;
   wire n_8_359;
   wire n_8_360;
   wire n_8_361;
   wire n_8_0_44;
   wire n_8_362;
   wire n_8_363;
   wire n_8_364;
   wire n_8_365;
   wire n_8_366;
   wire n_8_367;
   wire n_8_368;
   wire n_8_369;
   wire n_8_370;
   wire n_8_371;
   wire n_8_372;
   wire n_8_373;
   wire n_8_374;
   wire n_8_375;
   wire n_8_376;
   wire n_8_377;
   wire n_8_378;
   wire n_8_379;
   wire n_8_380;
   wire n_8_381;
   wire n_8_382;
   wire n_8_383;
   wire n_8_384;
   wire n_8_385;
   wire n_8_386;
   wire n_8_387;
   wire n_8_388;
   wire n_8_389;
   wire n_8_390;
   wire n_8_391;
   wire n_8_392;
   wire n_8_393;
   wire n_8_394;
   wire n_8_0_45;
   wire n_8_1026;
   wire n_8_1027;
   wire n_8_1028;
   wire n_8_1029;
   wire n_8_1030;
   wire n_8_1031;
   wire n_8_1032;
   wire n_8_1033;
   wire n_8_1034;
   wire n_8_1035;
   wire n_8_1036;
   wire n_8_1037;
   wire n_8_1038;
   wire n_8_1039;
   wire n_8_1040;
   wire n_8_1041;
   wire n_8_1042;
   wire n_8_1043;
   wire n_8_1044;
   wire n_8_1045;
   wire n_8_1046;
   wire n_8_1047;
   wire n_8_1048;
   wire n_8_1049;
   wire n_8_1050;
   wire n_8_1051;
   wire n_8_1052;
   wire n_8_1053;
   wire n_8_1054;
   wire n_8_395;
   wire n_8_396;
   wire n_8_397;
   wire n_8_398;
   wire n_8_0_46;
   wire n_8_981;
   wire n_8_982;
   wire n_8_983;
   wire n_8_984;
   wire n_8_985;
   wire n_8_986;
   wire n_8_987;
   wire n_8_988;
   wire n_8_989;
   wire n_8_990;
   wire n_8_991;
   wire n_8_992;
   wire n_8_993;
   wire n_8_994;
   wire n_8_995;
   wire n_8_996;
   wire n_8_997;
   wire n_8_998;
   wire n_8_999;
   wire n_8_1000;
   wire n_8_1001;
   wire n_8_1002;
   wire n_8_1003;
   wire n_8_1004;
   wire n_8_1005;
   wire n_8_1006;
   wire n_8_1007;
   wire n_8_1008;
   wire n_8_1009;
   wire n_8_1010;
   wire n_8_1011;
   wire n_8_1012;
   wire n_8_1024;
   wire n_8_0_47;
   wire n_8_935;
   wire n_8_936;
   wire n_8_937;
   wire n_8_938;
   wire n_8_939;
   wire n_8_940;
   wire n_8_941;
   wire n_8_942;
   wire n_8_943;
   wire n_8_944;
   wire n_8_945;
   wire n_8_946;
   wire n_8_947;
   wire n_8_948;
   wire n_8_949;
   wire n_8_950;
   wire n_8_951;
   wire n_8_952;
   wire n_8_953;
   wire n_8_954;
   wire n_8_955;
   wire n_8_956;
   wire n_8_957;
   wire n_8_958;
   wire n_8_959;
   wire n_8_960;
   wire n_8_961;
   wire n_8_962;
   wire n_8_963;
   wire n_8_964;
   wire n_8_965;
   wire n_8_966;
   wire n_8_979;
   wire n_8_0_48;
   wire n_8_888;
   wire n_8_889;
   wire n_8_890;
   wire n_8_891;
   wire n_8_892;
   wire n_8_893;
   wire n_8_894;
   wire n_8_895;
   wire n_8_896;
   wire n_8_897;
   wire n_8_898;
   wire n_8_899;
   wire n_8_900;
   wire n_8_901;
   wire n_8_902;
   wire n_8_903;
   wire n_8_904;
   wire n_8_905;
   wire n_8_906;
   wire n_8_907;
   wire n_8_908;
   wire n_8_909;
   wire n_8_910;
   wire n_8_911;
   wire n_8_912;
   wire n_8_913;
   wire n_8_914;
   wire n_8_915;
   wire n_8_916;
   wire n_8_917;
   wire n_8_918;
   wire n_8_919;
   wire n_8_933;
   wire n_8_0_49;
   wire n_8_840;
   wire n_8_841;
   wire n_8_842;
   wire n_8_843;
   wire n_8_844;
   wire n_8_845;
   wire n_8_846;
   wire n_8_847;
   wire n_8_848;
   wire n_8_849;
   wire n_8_850;
   wire n_8_851;
   wire n_8_852;
   wire n_8_853;
   wire n_8_854;
   wire n_8_855;
   wire n_8_856;
   wire n_8_857;
   wire n_8_858;
   wire n_8_859;
   wire n_8_860;
   wire n_8_861;
   wire n_8_862;
   wire n_8_863;
   wire n_8_864;
   wire n_8_865;
   wire n_8_866;
   wire n_8_867;
   wire n_8_868;
   wire n_8_869;
   wire n_8_870;
   wire n_8_871;
   wire n_8_886;
   wire n_8_0_50;
   wire n_8_791;
   wire n_8_792;
   wire n_8_793;
   wire n_8_794;
   wire n_8_795;
   wire n_8_796;
   wire n_8_797;
   wire n_8_798;
   wire n_8_799;
   wire n_8_800;
   wire n_8_801;
   wire n_8_802;
   wire n_8_803;
   wire n_8_804;
   wire n_8_805;
   wire n_8_806;
   wire n_8_807;
   wire n_8_808;
   wire n_8_809;
   wire n_8_810;
   wire n_8_811;
   wire n_8_812;
   wire n_8_813;
   wire n_8_814;
   wire n_8_815;
   wire n_8_816;
   wire n_8_817;
   wire n_8_818;
   wire n_8_819;
   wire n_8_820;
   wire n_8_821;
   wire n_8_822;
   wire n_8_838;
   wire n_8_0_51;
   wire n_8_741;
   wire n_8_742;
   wire n_8_743;
   wire n_8_744;
   wire n_8_745;
   wire n_8_746;
   wire n_8_747;
   wire n_8_748;
   wire n_8_749;
   wire n_8_750;
   wire n_8_751;
   wire n_8_752;
   wire n_8_753;
   wire n_8_754;
   wire n_8_755;
   wire n_8_756;
   wire n_8_757;
   wire n_8_758;
   wire n_8_759;
   wire n_8_760;
   wire n_8_761;
   wire n_8_762;
   wire n_8_763;
   wire n_8_764;
   wire n_8_765;
   wire n_8_766;
   wire n_8_767;
   wire n_8_768;
   wire n_8_769;
   wire n_8_770;
   wire n_8_771;
   wire n_8_772;
   wire n_8_789;
   wire n_8_0_52;
   wire n_8_690;
   wire n_8_691;
   wire n_8_692;
   wire n_8_693;
   wire n_8_694;
   wire n_8_695;
   wire n_8_696;
   wire n_8_697;
   wire n_8_698;
   wire n_8_699;
   wire n_8_700;
   wire n_8_701;
   wire n_8_702;
   wire n_8_703;
   wire n_8_704;
   wire n_8_705;
   wire n_8_706;
   wire n_8_707;
   wire n_8_708;
   wire n_8_709;
   wire n_8_710;
   wire n_8_711;
   wire n_8_712;
   wire n_8_713;
   wire n_8_714;
   wire n_8_715;
   wire n_8_716;
   wire n_8_717;
   wire n_8_718;
   wire n_8_719;
   wire n_8_720;
   wire n_8_721;
   wire n_8_739;
   wire n_8_0_53;
   wire n_8_638;
   wire n_8_639;
   wire n_8_640;
   wire n_8_641;
   wire n_8_642;
   wire n_8_643;
   wire n_8_644;
   wire n_8_645;
   wire n_8_646;
   wire n_8_647;
   wire n_8_648;
   wire n_8_649;
   wire n_8_650;
   wire n_8_651;
   wire n_8_652;
   wire n_8_653;
   wire n_8_654;
   wire n_8_655;
   wire n_8_656;
   wire n_8_657;
   wire n_8_658;
   wire n_8_659;
   wire n_8_660;
   wire n_8_661;
   wire n_8_662;
   wire n_8_663;
   wire n_8_664;
   wire n_8_665;
   wire n_8_666;
   wire n_8_667;
   wire n_8_668;
   wire n_8_669;
   wire n_8_688;
   wire n_8_0_54;
   wire n_8_585;
   wire n_8_586;
   wire n_8_587;
   wire n_8_588;
   wire n_8_589;
   wire n_8_590;
   wire n_8_591;
   wire n_8_592;
   wire n_8_593;
   wire n_8_594;
   wire n_8_595;
   wire n_8_596;
   wire n_8_597;
   wire n_8_598;
   wire n_8_599;
   wire n_8_600;
   wire n_8_601;
   wire n_8_602;
   wire n_8_603;
   wire n_8_604;
   wire n_8_605;
   wire n_8_606;
   wire n_8_607;
   wire n_8_608;
   wire n_8_609;
   wire n_8_610;
   wire n_8_611;
   wire n_8_612;
   wire n_8_613;
   wire n_8_614;
   wire n_8_615;
   wire n_8_616;
   wire n_8_636;
   wire n_8_0_55;
   wire n_8_531;
   wire n_8_532;
   wire n_8_533;
   wire n_8_534;
   wire n_8_535;
   wire n_8_536;
   wire n_8_537;
   wire n_8_538;
   wire n_8_539;
   wire n_8_540;
   wire n_8_541;
   wire n_8_542;
   wire n_8_543;
   wire n_8_544;
   wire n_8_545;
   wire n_8_546;
   wire n_8_547;
   wire n_8_548;
   wire n_8_549;
   wire n_8_550;
   wire n_8_551;
   wire n_8_552;
   wire n_8_553;
   wire n_8_554;
   wire n_8_555;
   wire n_8_556;
   wire n_8_557;
   wire n_8_558;
   wire n_8_559;
   wire n_8_560;
   wire n_8_561;
   wire n_8_562;
   wire n_8_583;
   wire n_8_476;
   wire n_8_477;
   wire n_8_478;
   wire n_8_479;
   wire n_8_480;
   wire n_8_481;
   wire n_8_482;
   wire n_8_483;
   wire n_8_484;
   wire n_8_485;
   wire n_8_486;
   wire n_8_487;
   wire n_8_488;
   wire n_8_489;
   wire n_8_490;
   wire n_8_491;
   wire n_8_492;
   wire n_8_493;
   wire n_8_494;
   wire n_8_495;
   wire n_8_496;
   wire n_8_497;
   wire n_8_498;
   wire n_8_499;
   wire n_8_500;
   wire n_8_501;
   wire n_8_502;
   wire n_8_503;
   wire n_8_504;
   wire n_8_506;
   wire n_8_507;
   wire n_8_526;
   wire n_8_420;
   wire n_8_421;
   wire n_8_422;
   wire n_8_423;
   wire n_8_424;
   wire n_8_425;
   wire n_8_426;
   wire n_8_427;
   wire n_8_428;
   wire n_8_429;
   wire n_8_430;
   wire n_8_431;
   wire n_8_432;
   wire n_8_433;
   wire n_8_434;
   wire n_8_435;
   wire n_8_436;
   wire n_8_437;
   wire n_8_438;
   wire n_8_439;
   wire n_8_440;
   wire n_8_441;
   wire n_8_442;
   wire n_8_443;
   wire n_8_444;
   wire n_8_445;
   wire n_8_446;
   wire n_8_447;
   wire n_8_449;
   wire n_8_451;
   wire n_8_471;
   wire n_8_399;
   wire n_8_400;
   wire n_8_401;
   wire n_8_402;
   wire n_8_403;
   wire n_8_404;
   wire n_8_405;
   wire n_8_406;
   wire n_8_407;
   wire n_8_408;
   wire n_8_409;
   wire n_8_410;
   wire n_8_411;
   wire n_8_412;
   wire n_8_413;
   wire n_8_414;
   wire n_8_415;
   wire n_8_416;
   wire n_8_417;
   wire n_8_418;
   wire n_8_419;
   wire n_8_452;
   wire n_8_453;
   wire n_8_454;
   wire n_8_455;
   wire n_8_456;
   wire n_8_457;
   wire n_8_458;
   wire n_8_459;
   wire n_8_461;
   wire n_8_463;
   wire n_8_464;
   wire n_8_465;
   wire n_8_466;
   wire n_8_467;
   wire n_8_468;
   wire n_8_469;
   wire n_8_470;
   wire n_8_472;
   wire n_8_473;
   wire n_8_474;
   wire n_8_475;
   wire n_8_508;
   wire n_8_509;
   wire n_8_510;
   wire n_8_511;
   wire n_8_512;
   wire n_8_513;
   wire n_8_514;
   wire n_8_515;
   wire n_8_516;
   wire n_8_517;
   wire n_8_518;
   wire n_8_519;
   wire n_8_520;
   wire n_8_521;
   wire n_8_522;
   wire n_8_523;
   wire n_8_524;
   wire n_8_525;
   wire n_8_529;
   wire n_8_563;
   wire n_8_564;
   wire n_8_565;
   wire n_8_566;
   wire n_8_567;
   wire n_8_568;
   wire n_8_569;
   wire n_8_570;
   wire n_8_571;
   wire n_8_572;
   wire n_8_573;
   wire n_8_574;
   wire n_8_575;
   wire n_8_576;
   wire n_8_577;
   wire n_8_578;
   wire n_8_579;
   wire n_8_580;
   wire n_8_581;
   wire n_8_582;
   wire n_8_584;
   wire n_8_617;
   wire n_8_618;
   wire n_8_619;
   wire n_8_620;
   wire n_8_621;
   wire n_8_622;
   wire n_8_623;
   wire n_8_624;
   wire n_8_625;
   wire n_8_626;
   wire n_8_629;
   wire n_8_630;
   wire n_8_631;
   wire n_8_632;
   wire n_8_633;
   wire n_8_634;
   wire n_8_635;
   wire n_8_637;
   wire n_8_670;
   wire n_8_671;
   wire n_8_672;
   wire n_8_673;
   wire n_8_674;
   wire n_8_675;
   wire n_8_676;
   wire n_8_677;
   wire n_8_678;
   wire n_8_679;
   wire n_8_680;
   wire n_8_681;
   wire n_8_682;
   wire n_8_683;
   wire n_8_684;
   wire n_8_685;
   wire n_8_687;
   wire n_8_689;
   wire n_8_722;
   wire n_8_723;
   wire n_8_725;
   wire n_8_726;
   wire n_8_728;
   wire n_8_729;
   wire n_8_730;
   wire n_8_731;
   wire n_8_732;
   wire n_8_733;
   wire n_8_734;
   wire n_8_735;
   wire n_8_736;
   wire n_8_737;
   wire n_8_738;
   wire n_8_740;
   wire n_8_773;
   wire n_8_774;
   wire n_8_775;
   wire n_8_776;
   wire n_8_777;
   wire n_8_778;
   wire n_8_779;
   wire n_8_780;
   wire n_8_781;
   wire n_8_782;
   wire n_8_783;
   wire n_8_784;
   wire n_8_785;
   wire n_8_787;
   wire n_8_788;
   wire n_8_790;
   wire n_8_824;
   wire n_8_825;
   wire n_8_826;
   wire n_8_827;
   wire n_8_828;
   wire n_8_829;
   wire n_8_830;
   wire n_8_831;
   wire n_8_832;
   wire n_8_833;
   wire n_8_834;
   wire n_8_835;
   wire n_8_836;
   wire n_8_837;
   wire n_8_839;
   wire n_8_872;
   wire n_8_873;
   wire n_8_874;
   wire n_8_875;
   wire n_8_876;
   wire n_8_877;
   wire n_8_878;
   wire n_8_879;
   wire n_8_880;
   wire n_8_881;
   wire n_8_882;
   wire n_8_883;
   wire n_8_884;
   wire n_8_885;
   wire n_8_920;
   wire n_8_922;
   wire n_8_923;
   wire n_8_924;
   wire n_8_925;
   wire n_8_926;
   wire n_8_927;
   wire n_8_928;
   wire n_8_929;
   wire n_8_930;
   wire n_8_931;
   wire n_8_932;
   wire n_8_934;
   wire n_8_967;
   wire n_8_968;
   wire n_8_969;
   wire n_8_970;
   wire n_8_971;
   wire n_8_972;
   wire n_8_973;
   wire n_8_974;
   wire n_8_975;
   wire n_8_976;
   wire n_8_977;
   wire n_8_978;
   wire n_8_980;
   wire n_8_1013;
   wire n_8_1014;
   wire n_8_1015;
   wire n_8_1016;
   wire n_8_1017;
   wire n_8_1018;
   wire n_8_1020;
   wire n_8_1022;
   wire n_8_1023;
   wire n_8_1025;
   wire n_8_0_65;
   wire n_8_0_66;
   wire n_8_0_67;
   wire n_8_0_68;
   wire n_8_0_69;
   wire n_8_0_70;
   wire n_8_0_71;
   wire n_8_0_72;
   wire n_8_0_73;
   wire n_8_0_74;
   wire n_8_0_75;
   wire n_8_0_76;
   wire n_8_0_77;
   wire n_8_0_78;
   wire n_8_0_79;
   wire n_8_0_80;
   wire n_8_0_81;
   wire n_8_0_82;
   wire n_8_0_83;
   wire n_8_0_84;
   wire n_8_0_85;
   wire n_8_0_86;
   wire n_8_0_87;
   wire n_8_0_88;
   wire n_8_0_89;
   wire n_8_0_90;
   wire n_8_0_91;
   wire n_8_0_92;
   wire n_8_0_93;
   wire n_8_0_94;
   wire n_8_0_95;
   wire n_8_0_96;
   wire n_8_0_97;
   wire n_8_25;
   wire n_8_27;
   wire n_8_28;
   wire n_8_65;
   wire n_8_98;
   wire n_8_99;
   wire n_8_100;
   wire n_8_131;
   wire n_8_133;
   wire n_8_164;
   wire n_8_197;
   wire n_8_198;
   wire n_8_199;
   wire n_8_231;
   wire n_8_232;
   wire n_8_233;
   wire n_8_234;
   wire n_8_236;
   wire n_8_238;
   wire n_8_240;
   wire n_8_241;
   wire n_8_242;
   wire n_8_505;
   wire n_8_448;
   wire n_8_450;
   wire n_8_460;
   wire n_8_462;
   wire n_8_527;
   wire n_8_528;
   wire n_8_530;
   wire n_8_627;
   wire n_8_628;
   wire n_8_686;
   wire n_8_724;
   wire n_8_786;
   wire n_8_823;
   wire n_8_887;
   wire n_8_921;
   wire n_8_1019;
   wire n_8_1021;
   wire n_8_0_64;
   wire n_8_0_63;
   wire n_8_0_62;
   wire n_8_0_61;
   wire n_8_0_60;
   wire n_8_0_59;
   wire n_8_0_58;
   wire n_8_0_57;
   wire n_8_0_56;
   wire n_8_0_40;
   wire n_8_0_39;
   wire n_8_0_38;
   wire n_8_0_37;
   wire n_8_0_36;
   wire n_8_0_35;
   wire n_8_0_33;
   wire n_8_0_32;
   wire n_8_0_31;
   wire n_8_0_30;
   wire n_8_0_29;
   wire n_8_0_28;
   wire n_8_0_27;
   wire n_8_0_26;
   wire n_8_0_25;
   wire n_8_0_13;
   wire n_8_0_12;
   wire n_8_0_11;
   wire n_8_0_9;
   wire n_8_0_7;
   wire n_8_0_5;
   wire n_8_0_4;
   wire n_8_0_3;
   wire n_8_0_2;
   wire n_8_0_1;
   wire n_8_0_0;
   wire n_8_0_98;
   wire n_8_0_99;
   wire n_8_727;
   wire n_8_0_100;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_0_0;
   wire n_1_0_1;
   wire n_1_0_2;
   wire n_1_0_3;
   wire n_1_0_4;
   wire n_1_0_5;
   wire n_1_0_6;
   wire n_1_0_7;
   wire n_1_0_8;
   wire n_1_0_9;
   wire n_1_0_10;
   wire n_1_0_11;
   wire n_1_0_12;
   wire n_1_0_13;
   wire n_1_0_14;
   wire n_1_0_15;
   wire n_1_0_16;
   wire n_1_0_17;
   wire n_1_0_18;
   wire n_1_0_19;
   wire n_1_0_20;
   wire n_1_0_21;
   wire n_1_0_22;
   wire n_1_0_23;
   wire n_1_0_24;
   wire n_1_0_25;
   wire n_1_0_26;
   wire n_1_0_27;
   wire n_1_0_28;
   wire n_1_0_29;
   wire n_1_0_30;
   wire n_1_0_31;
   wire n_1_0_32;
   wire n_1_0_33;
   wire n_1_0_34;
   wire n_1_0_35;
   wire n_1_0_36;
   wire n_1_0_37;
   wire n_1_0_38;
   wire n_1_0_39;
   wire n_1_0_40;
   wire n_1_0_41;
   wire n_1_0_42;
   wire n_1_0_43;
   wire n_1_0_44;
   wire n_1_0_45;
   wire n_1_0_46;
   wire n_1_0_47;
   wire n_1_0_48;
   wire n_1_0_49;
   wire n_1_0_50;
   wire n_1_0_51;
   wire n_1_0_52;
   wire n_1_0_53;
   wire n_1_0_54;
   wire n_1_0_55;
   wire n_1_0_56;
   wire n_1_0_57;
   wire n_1_0_58;
   wire n_1_0_59;
   wire n_1_0_60;
   wire n_1_0_61;
   wire n_1_0_62;
   wire n_1_0_63;
   wire n_1_0_64;
   wire n_1_0_65;
   wire n_1_0_66;
   wire n_1_0_67;
   wire n_1_0_68;
   wire n_1_0_69;
   wire n_1_0_70;
   wire n_1_0_71;
   wire n_1_0_72;
   wire n_1_0_73;
   wire n_1_0_74;
   wire n_1_0_75;
   wire n_1_0_76;
   wire n_1_0_77;
   wire n_1_0_78;
   wire n_1_0_79;
   wire n_1_0_80;
   wire n_1_0_81;
   wire n_1_0_82;
   wire n_1_0_83;
   wire n_1_0_84;
   wire n_1_0_85;
   wire n_1_0_86;
   wire n_1_0_87;
   wire n_1_0_88;
   wire n_1_0_89;
   wire n_1_0_90;
   wire n_1_0_91;
   wire n_1_0_92;
   wire n_1_0_93;
   wire n_1_0_94;
   wire n_1_0_95;
   wire n_1_0_96;
   wire n_1_0_97;
   wire n_1_0_98;
   wire n_1_0_99;
   wire n_1_0_100;
   wire n_1_0_101;

   datapath__0_130 i_8_32 (.p_0({uc_0, uc_1, uc_2, uc_3, n_8_1025, uc_4, uc_5, 
      uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, 
      uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, 
      uc_27, uc_28, uc_29, n_8_1023, n_8_1022, n_8_1021, n_8_1020, n_8_1019, 
      n_8_1018, n_8_1017, n_8_1016, n_8_1015, n_8_1014, n_8_1013, n_8_980, 
      n_8_978, n_8_977, n_8_976, n_8_975, n_8_974, n_8_973, n_8_972, n_8_971, 
      n_8_970, n_8_969, n_8_968, n_8_967, n_8_934, n_8_932, n_8_931, n_8_930, 
      n_8_929, n_8_928, n_8_927, n_8_926, uc_30}), .p_1({uc_31, uc_32, uc_33, 
      uc_34, n_8_925, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, 
      uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, n_8_924, n_8_923, n_8_922, 
      n_8_921, n_8_920, n_8_887, n_8_885, n_8_884, n_8_883, n_8_882, n_8_881, 
      n_8_880, n_8_879, n_8_878, n_8_877, n_8_876, n_8_875, n_8_874, n_8_873, 
      n_8_872, n_8_839, n_8_837, n_8_836, n_8_835, n_8_834, n_8_833, n_8_832, 
      n_8_831, n_8_830, n_8_829, n_8_828, n_8_827, uc_60, uc_61}), .p_2({uc_62, 
      uc_63, uc_64, uc_65, n_8_826, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, 
      uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, 
      uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, n_8_825, n_8_824, 
      n_8_823, n_8_790, n_8_788, n_8_787, n_8_786, n_8_785, n_8_784, n_8_783, 
      n_8_782, n_8_781, n_8_780, n_8_779, n_8_778, n_8_777, n_8_776, n_8_775, 
      n_8_774, n_8_773, n_8_740, n_8_738, n_8_737, n_8_736, n_8_735, n_8_734, 
      n_8_733, n_8_732, n_8_731, n_8_730, n_8_729, n_8_728, uc_90, uc_91, uc_92}), 
      .p_3({uc_93, uc_94, uc_95, uc_96, n_8_727, uc_97, uc_98, uc_99, uc_100, 
      uc_101, uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, 
      uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, 
      uc_119, n_8_726, n_8_725, n_8_724, n_8_723, n_8_722, n_8_689, n_8_687, 
      n_8_686, n_8_685, n_8_684, n_8_683, n_8_682, n_8_681, n_8_680, n_8_679, 
      n_8_678, n_8_677, n_8_676, n_8_675, n_8_674, n_8_673, n_8_672, n_8_671, 
      n_8_670, n_8_637, n_8_635, n_8_634, n_8_633, n_8_632, n_8_631, n_8_630, 
      n_8_629, uc_120, uc_121, uc_122, uc_123}), .p_4({uc_124, uc_125, uc_126, 
      uc_127, n_8_628, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, 
      uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, 
      uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, n_8_627, n_8_626, n_8_625, 
      n_8_624, n_8_623, n_8_622, n_8_621, n_8_620, n_8_619, n_8_618, n_8_617, 
      n_8_584, n_8_582, n_8_581, n_8_580, n_8_579, n_8_578, n_8_577, n_8_576, 
      n_8_575, n_8_574, n_8_573, n_8_572, n_8_571, n_8_570, n_8_569, n_8_568, 
      n_8_567, n_8_566, n_8_565, n_8_564, n_8_563, uc_150, uc_151, uc_152, 
      uc_153, uc_154}), .p_5({uc_155, uc_156, uc_157, uc_158, n_8_530, uc_159, 
      uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, uc_168, 
      uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, uc_177, 
      uc_178, uc_179, n_8_529, n_8_528, n_8_527, n_8_525, n_8_524, n_8_523, 
      n_8_522, n_8_521, n_8_520, n_8_519, n_8_518, n_8_517, n_8_516, n_8_515, 
      n_8_514, n_8_513, n_8_512, n_8_511, n_8_510, n_8_509, n_8_508, n_8_475, 
      n_8_474, n_8_473, n_8_472, n_8_470, n_8_469, n_8_468, n_8_467, n_8_466, 
      n_8_465, n_8_464, uc_180, uc_181, uc_182, uc_183, uc_184, uc_185}), 
      .p_6({uc_186, uc_187, uc_188, uc_189, n_8_463, uc_190, uc_191, uc_192, 
      uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, 
      uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, uc_209, n_8_462, 
      n_8_461, n_8_460, n_8_459, n_8_458, n_8_457, n_8_456, n_8_455, n_8_454, 
      n_8_453, n_8_452, n_8_419, n_8_418, n_8_417, n_8_416, n_8_415, n_8_414, 
      n_8_413, n_8_412, n_8_411, n_8_410, n_8_409, n_8_408, n_8_407, n_8_406, 
      n_8_405, n_8_404, n_8_403, n_8_402, n_8_401, n_8_400, n_8_399, uc_210, 
      uc_211, uc_212, uc_213, uc_214, uc_215, uc_216}), .p_7({uc_217, uc_218, 
      uc_219, uc_220, n_8_471, uc_221, uc_222, uc_223, uc_224, uc_225, uc_226, 
      uc_227, uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, uc_234, uc_235, 
      uc_236, uc_237, uc_238, uc_239, n_8_451, n_8_450, n_8_449, n_8_448, 
      n_8_447, n_8_446, n_8_445, n_8_444, n_8_443, n_8_442, n_8_441, n_8_440, 
      n_8_439, n_8_438, n_8_437, n_8_436, n_8_435, n_8_434, n_8_433, n_8_432, 
      n_8_431, n_8_430, n_8_429, n_8_428, n_8_427, n_8_426, n_8_425, n_8_424, 
      n_8_423, n_8_422, n_8_421, n_8_420, uc_240, uc_241, uc_242, uc_243, uc_244, 
      uc_245, uc_246, uc_247}), .p_8({uc_248, uc_249, uc_250, uc_251, n_8_526, 
      uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, 
      uc_261, uc_262, uc_263, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, 
      n_8_507, n_8_506, n_8_505, n_8_504, n_8_503, n_8_502, n_8_501, n_8_500, 
      n_8_499, n_8_498, n_8_497, n_8_496, n_8_495, n_8_494, n_8_493, n_8_492, 
      n_8_491, n_8_490, n_8_489, n_8_488, n_8_487, n_8_486, n_8_485, n_8_484, 
      n_8_483, n_8_482, n_8_481, n_8_480, n_8_479, n_8_478, n_8_477, n_8_476, 
      uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, uc_278}), 
      .p_9({uc_279, n_8_583, uc_280, uc_281, uc_282, uc_283, uc_284, uc_285, 
      uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, 
      uc_295, uc_296, uc_297, uc_298, uc_299, n_8_562, n_8_561, n_8_560, n_8_559, 
      n_8_558, n_8_557, n_8_556, n_8_555, n_8_554, n_8_553, n_8_552, n_8_551, 
      n_8_550, n_8_549, n_8_548, n_8_547, n_8_546, n_8_545, n_8_544, n_8_543, 
      n_8_542, n_8_541, n_8_540, n_8_539, n_8_538, n_8_537, n_8_536, n_8_535, 
      n_8_534, n_8_533, n_8_532, n_8_531, uc_300, uc_301, uc_302, uc_303, uc_304, 
      uc_305, uc_306, uc_307, uc_308, uc_309}), .p_10({uc_310, n_8_636, uc_311, 
      uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, uc_319, uc_320, 
      uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, 
      n_8_616, n_8_615, n_8_614, n_8_613, n_8_612, n_8_611, n_8_610, n_8_609, 
      n_8_608, n_8_607, n_8_606, n_8_605, n_8_604, n_8_603, n_8_602, n_8_601, 
      n_8_600, n_8_599, n_8_598, n_8_597, n_8_596, n_8_595, n_8_594, n_8_593, 
      n_8_592, n_8_591, n_8_590, n_8_589, n_8_588, n_8_587, n_8_586, n_8_585, 
      uc_330, uc_331, uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, uc_338, 
      uc_339, uc_340}), .p_11({uc_341, n_8_688, uc_342, uc_343, uc_344, uc_345, 
      uc_346, uc_347, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, 
      uc_355, uc_356, uc_357, uc_358, uc_359, n_8_669, n_8_668, n_8_667, n_8_666, 
      n_8_665, n_8_664, n_8_663, n_8_662, n_8_661, n_8_660, n_8_659, n_8_658, 
      n_8_657, n_8_656, n_8_655, n_8_654, n_8_653, n_8_652, n_8_651, n_8_650, 
      n_8_649, n_8_648, n_8_647, n_8_646, n_8_645, n_8_644, n_8_643, n_8_642, 
      n_8_641, n_8_640, n_8_639, n_8_638, uc_360, uc_361, uc_362, uc_363, uc_364, 
      uc_365, uc_366, uc_367, uc_368, uc_369, uc_370, uc_371}), .p_12({uc_372, 
      n_8_739, uc_373, uc_374, uc_375, uc_376, uc_377, uc_378, uc_379, uc_380, 
      uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, 
      n_8_721, n_8_720, n_8_719, n_8_718, n_8_717, n_8_716, n_8_715, n_8_714, 
      n_8_713, n_8_712, n_8_711, n_8_710, n_8_709, n_8_708, n_8_707, n_8_706, 
      n_8_705, n_8_704, n_8_703, n_8_702, n_8_701, n_8_700, n_8_699, n_8_698, 
      n_8_697, n_8_696, n_8_695, n_8_694, n_8_693, n_8_692, n_8_691, n_8_690, 
      uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, 
      uc_399, uc_400, uc_401, uc_402}), .p_13({uc_403, n_8_789, uc_404, uc_405, 
      uc_406, uc_407, uc_408, uc_409, uc_410, uc_411, uc_412, uc_413, uc_414, 
      uc_415, uc_416, uc_417, uc_418, uc_419, n_8_772, n_8_771, n_8_770, n_8_769, 
      n_8_768, n_8_767, n_8_766, n_8_765, n_8_764, n_8_763, n_8_762, n_8_761, 
      n_8_760, n_8_759, n_8_758, n_8_757, n_8_756, n_8_755, n_8_754, n_8_753, 
      n_8_752, n_8_751, n_8_750, n_8_749, n_8_748, n_8_747, n_8_746, n_8_745, 
      n_8_744, n_8_743, n_8_742, n_8_741, uc_420, uc_421, uc_422, uc_423, uc_424, 
      uc_425, uc_426, uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, uc_433}), 
      .p_14({uc_434, n_8_838, uc_435, uc_436, uc_437, uc_438, uc_439, uc_440, 
      uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, 
      n_8_822, n_8_821, n_8_820, n_8_819, n_8_818, n_8_817, n_8_816, n_8_815, 
      n_8_814, n_8_813, n_8_812, n_8_811, n_8_810, n_8_809, n_8_808, n_8_807, 
      n_8_806, n_8_805, n_8_804, n_8_803, n_8_802, n_8_801, n_8_800, n_8_799, 
      n_8_798, n_8_797, n_8_796, n_8_795, n_8_794, n_8_793, n_8_792, n_8_791, 
      uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, 
      uc_459, uc_460, uc_461, uc_462, uc_463, uc_464}), .p_15({uc_465, n_8_886, 
      uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, uc_474, 
      uc_475, uc_476, uc_477, uc_478, uc_479, n_8_871, n_8_870, n_8_869, n_8_868, 
      n_8_867, n_8_866, n_8_865, n_8_864, n_8_863, n_8_862, n_8_861, n_8_860, 
      n_8_859, n_8_858, n_8_857, n_8_856, n_8_855, n_8_854, n_8_853, n_8_852, 
      n_8_851, n_8_850, n_8_849, n_8_848, n_8_847, n_8_846, n_8_845, n_8_844, 
      n_8_843, n_8_842, n_8_841, n_8_840, uc_480, uc_481, uc_482, uc_483, uc_484, 
      uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, uc_492, uc_493, 
      uc_494, uc_495}), .p_16({uc_496, n_8_933, uc_497, uc_498, uc_499, uc_500, 
      uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, 
      n_8_919, n_8_918, n_8_917, n_8_916, n_8_915, n_8_914, n_8_913, n_8_912, 
      n_8_911, n_8_910, n_8_909, n_8_908, n_8_907, n_8_906, n_8_905, n_8_904, 
      n_8_903, n_8_902, n_8_901, n_8_900, n_8_899, n_8_898, n_8_897, n_8_896, 
      n_8_895, n_8_894, n_8_893, n_8_892, n_8_891, n_8_890, n_8_889, n_8_888, 
      uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, uc_517, uc_518, 
      uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, uc_526}), .p_17({
      uc_527, n_8_979, uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, 
      uc_535, uc_536, uc_537, uc_538, uc_539, n_8_966, n_8_965, n_8_964, n_8_963, 
      n_8_962, n_8_961, n_8_960, n_8_959, n_8_958, n_8_957, n_8_956, n_8_955, 
      n_8_954, n_8_953, n_8_952, n_8_951, n_8_950, n_8_949, n_8_948, n_8_947, 
      n_8_946, n_8_945, n_8_944, n_8_943, n_8_942, n_8_941, n_8_940, n_8_939, 
      n_8_938, n_8_937, n_8_936, n_8_935, uc_540, uc_541, uc_542, uc_543, uc_544, 
      uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, 
      uc_554, uc_555, uc_556, uc_557}), .p_18({uc_558, n_8_1024, uc_559, uc_560, 
      uc_561, uc_562, uc_563, uc_564, uc_565, uc_566, uc_567, uc_568, uc_569, 
      n_8_1012, n_8_1011, n_8_1010, n_8_1009, n_8_1008, n_8_1007, n_8_1006, 
      n_8_1005, n_8_1004, n_8_1003, n_8_1002, n_8_1001, n_8_1000, n_8_999, 
      n_8_998, n_8_997, n_8_996, n_8_995, n_8_994, n_8_993, n_8_992, n_8_991, 
      n_8_990, n_8_989, n_8_988, n_8_987, n_8_986, n_8_985, n_8_984, n_8_983, 
      n_8_982, n_8_981, uc_570, uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, 
      uc_577, uc_578, uc_579, uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, 
      uc_586, uc_587, uc_588}), .p_19({uc_589, n_8_398, uc_590, uc_591, uc_592, 
      uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, n_8_397, n_8_396, 
      n_8_395, n_8_1054, n_8_1053, n_8_1052, n_8_1051, n_8_1050, n_8_1049, 
      n_8_1048, n_8_1047, n_8_1046, n_8_1045, n_8_1044, n_8_1043, n_8_1042, 
      n_8_1041, n_8_1040, n_8_1039, n_8_1038, n_8_1037, n_8_1036, n_8_1035, 
      n_8_1034, n_8_1033, n_8_1032, n_8_1031, n_8_1030, n_8_1029, n_8_1028, 
      n_8_1027, n_8_1026, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, 
      uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, 
      uc_616, uc_617, uc_618, uc_619}), .p_20({uc_620, n_8_394, uc_621, uc_622, 
      uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, uc_629, n_8_393, n_8_392, 
      n_8_391, n_8_390, n_8_389, n_8_388, n_8_387, n_8_386, n_8_385, n_8_384, 
      n_8_383, n_8_382, n_8_381, n_8_380, n_8_379, n_8_378, n_8_377, n_8_376, 
      n_8_375, n_8_374, n_8_373, n_8_372, n_8_371, n_8_370, n_8_369, n_8_368, 
      n_8_367, n_8_366, n_8_365, n_8_364, n_8_363, n_8_362, uc_630, uc_631, 
      uc_632, uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639, uc_640, 
      uc_641, uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, 
      uc_650}), .p_21({uc_651, n_8_361, uc_652, uc_653, uc_654, uc_655, uc_656, 
      uc_657, uc_658, uc_659, n_8_360, n_8_359, n_8_358, n_8_357, n_8_356, 
      n_8_355, n_8_354, n_8_353, n_8_352, n_8_351, n_8_350, n_8_349, n_8_348, 
      n_8_347, n_8_346, n_8_345, n_8_344, n_8_343, n_8_342, n_8_341, n_8_340, 
      n_8_339, n_8_338, n_8_337, n_8_336, n_8_335, n_8_334, n_8_333, n_8_332, 
      n_8_331, n_8_330, n_8_329, uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, 
      uc_666, uc_667, uc_668, uc_669, uc_670, uc_671, uc_672, uc_673, uc_674, 
      uc_675, uc_676, uc_677, uc_678, uc_679, uc_680, uc_681}), .p_22({uc_682, 
      n_8_328, uc_683, uc_684, uc_685, uc_686, uc_687, uc_688, uc_689, n_8_327, 
      n_8_326, n_8_325, n_8_324, n_8_323, n_8_322, n_8_321, n_8_320, n_8_319, 
      n_8_318, n_8_317, n_8_316, n_8_315, n_8_314, n_8_313, n_8_312, n_8_311, 
      n_8_310, n_8_309, n_8_308, n_8_307, n_8_306, n_8_305, n_8_304, n_8_303, 
      n_8_302, n_8_301, n_8_300, n_8_299, n_8_298, n_8_297, n_8_296, uc_690, 
      uc_691, uc_692, uc_693, uc_694, uc_695, uc_696, uc_697, uc_698, uc_699, 
      uc_700, uc_701, uc_702, uc_703, uc_704, uc_705, uc_706, uc_707, uc_708, 
      uc_709, uc_710, uc_711, uc_712}), .p_23({uc_713, n_8_295, uc_714, uc_715, 
      uc_716, uc_717, uc_718, uc_719, n_8_294, n_8_293, n_8_292, n_8_291, 
      n_8_290, n_8_289, n_8_288, n_8_287, n_8_286, n_8_285, n_8_284, n_8_283, 
      n_8_282, n_8_281, n_8_280, n_8_279, n_8_278, n_8_277, n_8_276, n_8_275, 
      n_8_274, n_8_273, n_8_272, n_8_271, n_8_270, n_8_269, n_8_268, n_8_267, 
      n_8_266, n_8_265, n_8_264, n_8_263, uc_720, uc_721, uc_722, uc_723, uc_724, 
      uc_725, uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, 
      uc_734, uc_735, uc_736, uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, 
      uc_743}), .p_24({uc_744, n_8_262, uc_745, uc_746, uc_747, uc_748, uc_749, 
      n_8_261, n_8_260, n_8_259, n_8_258, n_8_257, n_8_256, n_8_255, n_8_254, 
      n_8_253, n_8_252, n_8_251, n_8_250, n_8_249, n_8_248, n_8_247, n_8_246, 
      n_8_245, n_8_244, n_8_243, n_8_242, n_8_241, n_8_240, n_8_239, n_8_238, 
      n_8_237, n_8_236, n_8_235, n_8_234, n_8_233, n_8_232, n_8_231, n_8_230, 
      uc_750, uc_751, uc_752, uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, 
      uc_759, uc_760, uc_761, uc_762, uc_763, uc_764, uc_765, uc_766, uc_767, 
      uc_768, uc_769, uc_770, uc_771, uc_772, uc_773, uc_774}), .p_25({uc_775, 
      n_8_229, uc_776, uc_777, uc_778, uc_779, n_8_228, n_8_227, n_8_226, 
      n_8_225, n_8_224, n_8_223, n_8_222, n_8_221, n_8_220, n_8_219, n_8_218, 
      n_8_217, n_8_216, n_8_215, n_8_214, n_8_213, n_8_212, n_8_211, n_8_210, 
      n_8_209, n_8_208, n_8_207, n_8_206, n_8_205, n_8_204, n_8_203, n_8_202, 
      n_8_201, n_8_200, n_8_199, n_8_198, n_8_197, uc_780, uc_781, uc_782, 
      uc_783, uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, 
      uc_792, uc_793, uc_794, uc_795, uc_796, uc_797, uc_798, uc_799, uc_800, 
      uc_801, uc_802, uc_803, uc_804, uc_805}), .p_26({uc_806, n_8_196, uc_807, 
      uc_808, uc_809, n_8_195, n_8_194, n_8_193, n_8_192, n_8_191, n_8_190, 
      n_8_189, n_8_188, n_8_187, n_8_186, n_8_185, n_8_184, n_8_183, n_8_182, 
      n_8_181, n_8_180, n_8_179, n_8_178, n_8_177, n_8_176, n_8_175, n_8_174, 
      n_8_173, n_8_172, n_8_171, n_8_170, n_8_169, n_8_168, n_8_167, n_8_166, 
      n_8_165, n_8_164, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, 
      uc_817, uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, 
      uc_826, uc_827, uc_828, uc_829, uc_830, uc_831, uc_832, uc_833, uc_834, 
      uc_835, uc_836}), .p_27({uc_837, uc_838, uc_839, n_8_163, n_8_162, n_8_161, 
      n_8_160, n_8_159, n_8_158, n_8_157, n_8_156, n_8_155, n_8_154, n_8_153, 
      n_8_152, n_8_151, n_8_150, n_8_149, n_8_148, n_8_147, n_8_146, n_8_145, 
      n_8_144, n_8_143, n_8_142, n_8_141, n_8_140, n_8_139, n_8_138, n_8_137, 
      n_8_136, n_8_135, n_8_134, n_8_133, n_8_132, n_8_131, uc_840, uc_841, 
      uc_842, uc_843, uc_844, uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, 
      uc_851, uc_852, uc_853, uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, 
      uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, uc_866, uc_867}), .p_28({
      uc_868, uc_869, n_8_130, n_8_129, n_8_128, n_8_127, n_8_126, n_8_125, 
      n_8_124, n_8_123, n_8_122, n_8_121, n_8_120, n_8_119, n_8_118, n_8_117, 
      n_8_116, n_8_115, n_8_114, n_8_113, n_8_112, n_8_111, n_8_110, n_8_109, 
      n_8_108, n_8_107, n_8_106, n_8_105, n_8_104, n_8_103, n_8_102, n_8_101, 
      n_8_100, n_8_99, n_8_98, uc_870, uc_871, uc_872, uc_873, uc_874, uc_875, 
      uc_876, uc_877, uc_878, uc_879, uc_880, uc_881, uc_882, uc_883, uc_884, 
      uc_885, uc_886, uc_887, uc_888, uc_889, uc_890, uc_891, uc_892, uc_893, 
      uc_894, uc_895, uc_896, uc_897, uc_898}), .p_29({uc_899, n_8_97, n_8_96, 
      n_8_95, n_8_94, n_8_93, n_8_92, n_8_91, n_8_90, n_8_89, n_8_88, n_8_87, 
      n_8_86, n_8_85, n_8_84, n_8_83, n_8_82, n_8_81, n_8_80, n_8_79, n_8_78, 
      n_8_77, n_8_76, n_8_75, n_8_74, n_8_73, n_8_72, n_8_71, n_8_70, n_8_69, 
      n_8_68, n_8_67, n_8_66, n_8_65, uc_900, uc_901, uc_902, uc_903, uc_904, 
      uc_905, uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, uc_912, uc_913, 
      uc_914, uc_915, uc_916, uc_917, uc_918, uc_919, uc_920, uc_921, uc_922, 
      uc_923, uc_924, uc_925, uc_926, uc_927, uc_928, uc_929}), .p_30({n_8_64, 
      n_8_63, n_8_62, n_8_61, n_8_60, n_8_59, n_8_58, n_8_57, n_8_56, n_8_55, 
      n_8_54, n_8_53, n_8_52, n_8_51, n_8_50, n_8_49, n_8_48, n_8_47, n_8_46, 
      n_8_45, n_8_44, n_8_43, n_8_42, n_8_41, n_8_40, n_8_39, n_8_38, n_8_37, 
      n_8_36, n_8_35, n_8_34, n_8_33, n_8_32, uc_930, uc_931, uc_932, uc_933, 
      uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, uc_940, uc_941, uc_942, 
      uc_943, uc_944, uc_945, uc_946, uc_947, uc_948, uc_949, uc_950, uc_951, 
      uc_952, uc_953, uc_954, uc_955, uc_956, uc_957, uc_958, uc_959, uc_960}), 
      .out({uc_961, uc_962, n_8_31, uc_963, uc_964, uc_965, uc_966, uc_967, 
      uc_968, uc_969, uc_970, uc_971, uc_972, uc_973, uc_974, uc_975, uc_976, 
      uc_977, uc_978, uc_979, uc_980, uc_981, uc_982, uc_983, uc_984, uc_985, 
      uc_986, uc_987, uc_988, uc_989, uc_990, uc_991, n_8_30, n_8_29, n_8_28, 
      n_8_27, n_8_26, n_8_25, n_8_24, n_8_23, n_8_22, n_8_21, n_8_20, n_8_19, 
      n_8_18, n_8_17, n_8_16, n_8_15, n_8_14, n_8_13, n_8_12, n_8_11, n_8_10, 
      n_8_9, n_8_8, n_8_7, n_8_6, n_8_5, n_8_4, n_8_3, n_8_2, n_8_1, n_8_0, 
      uc_992}), .out31({n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
      n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
      n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
      n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
      n_4, n_3, n_2, n_1, n_0, uc_993}));
   NOR2_X1 i_8_0_2 (.A1(n_8_0_0), .A2(n_8_0_1), .ZN(n_63));
   NOR2_X1 i_8_0_4 (.A1(n_8_0_0), .A2(n_8_0_2), .ZN(n_8_0));
   NOR2_X1 i_8_0_6 (.A1(n_8_0_0), .A2(n_8_0_3), .ZN(n_8_1));
   NOR2_X1 i_8_0_8 (.A1(n_8_0_0), .A2(n_8_0_4), .ZN(n_8_2));
   NOR2_X1 i_8_0_10 (.A1(n_8_0_0), .A2(n_8_0_5), .ZN(n_8_3));
   INV_X1 i_8_0_11 (.A(n_108), .ZN(n_8_0_6));
   NOR2_X1 i_8_0_12 (.A1(n_8_0_0), .A2(n_8_0_6), .ZN(n_8_4));
   NOR2_X1 i_8_0_14 (.A1(n_8_0_0), .A2(n_8_0_7), .ZN(n_8_5));
   INV_X1 i_8_0_15 (.A(n_110), .ZN(n_8_0_8));
   NOR2_X1 i_8_0_16 (.A1(n_8_0_0), .A2(n_8_0_8), .ZN(n_8_6));
   NOR2_X1 i_8_0_18 (.A1(n_8_0_0), .A2(n_8_0_9), .ZN(n_8_7));
   INV_X1 i_8_0_19 (.A(n_111), .ZN(n_8_0_10));
   NOR2_X1 i_8_0_20 (.A1(n_8_0_0), .A2(n_8_0_10), .ZN(n_8_8));
   NOR2_X1 i_8_0_22 (.A1(n_8_0_0), .A2(n_8_0_11), .ZN(n_8_9));
   NOR2_X1 i_8_0_24 (.A1(n_8_0_0), .A2(n_8_0_12), .ZN(n_8_10));
   NOR2_X1 i_8_0_26 (.A1(n_8_0_0), .A2(n_8_0_13), .ZN(n_8_11));
   INV_X1 i_8_0_27 (.A(n_115), .ZN(n_8_0_14));
   NOR2_X1 i_8_0_28 (.A1(n_8_0_0), .A2(n_8_0_14), .ZN(n_8_12));
   INV_X1 i_8_0_29 (.A(n_116), .ZN(n_8_0_15));
   NOR2_X1 i_8_0_30 (.A1(n_8_0_0), .A2(n_8_0_15), .ZN(n_8_13));
   INV_X1 i_8_0_31 (.A(n_126), .ZN(n_8_0_16));
   NOR2_X1 i_8_0_32 (.A1(n_8_0_0), .A2(n_8_0_16), .ZN(n_8_14));
   INV_X1 i_8_0_33 (.A(n_117), .ZN(n_8_0_17));
   NOR2_X1 i_8_0_34 (.A1(n_8_0_0), .A2(n_8_0_17), .ZN(n_8_15));
   INV_X1 i_8_0_35 (.A(n_118), .ZN(n_8_0_18));
   NOR2_X1 i_8_0_36 (.A1(n_8_0_0), .A2(n_8_0_18), .ZN(n_8_16));
   INV_X1 i_8_0_37 (.A(n_82), .ZN(n_8_0_19));
   NOR2_X1 i_8_0_38 (.A1(n_8_0_0), .A2(n_8_0_19), .ZN(n_8_17));
   INV_X1 i_8_0_39 (.A(n_119), .ZN(n_8_0_20));
   NOR2_X1 i_8_0_40 (.A1(n_8_0_0), .A2(n_8_0_20), .ZN(n_8_18));
   INV_X1 i_8_0_41 (.A(n_120), .ZN(n_8_0_21));
   NOR2_X1 i_8_0_42 (.A1(n_8_0_0), .A2(n_8_0_21), .ZN(n_8_19));
   INV_X1 i_8_0_43 (.A(n_83), .ZN(n_8_0_22));
   NOR2_X1 i_8_0_44 (.A1(n_8_0_0), .A2(n_8_0_22), .ZN(n_8_20));
   INV_X1 i_8_0_45 (.A(n_121), .ZN(n_8_0_23));
   NOR2_X1 i_8_0_46 (.A1(n_8_0_0), .A2(n_8_0_23), .ZN(n_8_21));
   INV_X1 i_8_0_47 (.A(n_72), .ZN(n_8_0_24));
   NOR2_X1 i_8_0_48 (.A1(n_8_0_0), .A2(n_8_0_24), .ZN(n_8_22));
   NOR2_X1 i_8_0_50 (.A1(n_8_0_0), .A2(n_8_0_25), .ZN(n_8_23));
   NOR2_X1 i_8_0_52 (.A1(n_8_0_0), .A2(n_8_0_26), .ZN(n_8_24));
   NOR2_X1 i_8_0_56 (.A1(n_8_0_0), .A2(n_8_0_28), .ZN(n_8_26));
   NOR2_X1 i_8_0_62 (.A1(n_8_0_0), .A2(n_8_0_31), .ZN(n_8_29));
   NOR2_X1 i_8_0_64 (.A1(n_8_0_0), .A2(n_8_0_32), .ZN(n_8_30));
   NOR2_X1 i_8_0_66 (.A1(n_8_0_0), .A2(n_8_0_33), .ZN(n_8_31));
   INV_X1 i_8_0_67 (.A(n_68), .ZN(n_8_0_34));
   NOR2_X1 i_8_0_68 (.A1(n_8_0_34), .A2(n_8_0_1), .ZN(n_8_32));
   NOR2_X1 i_8_0_69 (.A1(n_8_0_34), .A2(n_8_0_2), .ZN(n_8_33));
   NOR2_X1 i_8_0_70 (.A1(n_8_0_34), .A2(n_8_0_3), .ZN(n_8_34));
   NOR2_X1 i_8_0_71 (.A1(n_8_0_34), .A2(n_8_0_4), .ZN(n_8_35));
   NOR2_X1 i_8_0_72 (.A1(n_8_0_34), .A2(n_8_0_5), .ZN(n_8_36));
   NOR2_X1 i_8_0_73 (.A1(n_8_0_34), .A2(n_8_0_6), .ZN(n_8_37));
   NOR2_X1 i_8_0_74 (.A1(n_8_0_34), .A2(n_8_0_7), .ZN(n_8_38));
   NOR2_X1 i_8_0_75 (.A1(n_8_0_34), .A2(n_8_0_8), .ZN(n_8_39));
   NOR2_X1 i_8_0_76 (.A1(n_8_0_34), .A2(n_8_0_9), .ZN(n_8_40));
   NOR2_X1 i_8_0_77 (.A1(n_8_0_34), .A2(n_8_0_10), .ZN(n_8_41));
   NOR2_X1 i_8_0_78 (.A1(n_8_0_34), .A2(n_8_0_11), .ZN(n_8_42));
   NOR2_X1 i_8_0_79 (.A1(n_8_0_34), .A2(n_8_0_12), .ZN(n_8_43));
   NOR2_X1 i_8_0_80 (.A1(n_8_0_34), .A2(n_8_0_13), .ZN(n_8_44));
   NOR2_X1 i_8_0_81 (.A1(n_8_0_34), .A2(n_8_0_14), .ZN(n_8_45));
   NOR2_X1 i_8_0_82 (.A1(n_8_0_34), .A2(n_8_0_15), .ZN(n_8_46));
   NOR2_X1 i_8_0_83 (.A1(n_8_0_34), .A2(n_8_0_16), .ZN(n_8_47));
   NOR2_X1 i_8_0_84 (.A1(n_8_0_34), .A2(n_8_0_17), .ZN(n_8_48));
   NOR2_X1 i_8_0_85 (.A1(n_8_0_34), .A2(n_8_0_18), .ZN(n_8_49));
   NOR2_X1 i_8_0_86 (.A1(n_8_0_34), .A2(n_8_0_19), .ZN(n_8_50));
   NOR2_X1 i_8_0_87 (.A1(n_8_0_34), .A2(n_8_0_20), .ZN(n_8_51));
   NOR2_X1 i_8_0_88 (.A1(n_8_0_34), .A2(n_8_0_21), .ZN(n_8_52));
   NOR2_X1 i_8_0_89 (.A1(n_8_0_34), .A2(n_8_0_22), .ZN(n_8_53));
   NOR2_X1 i_8_0_90 (.A1(n_8_0_34), .A2(n_8_0_23), .ZN(n_8_54));
   NOR2_X1 i_8_0_91 (.A1(n_8_0_34), .A2(n_8_0_24), .ZN(n_8_55));
   NOR2_X1 i_8_0_92 (.A1(n_8_0_34), .A2(n_8_0_25), .ZN(n_8_56));
   NOR2_X1 i_8_0_93 (.A1(n_8_0_34), .A2(n_8_0_26), .ZN(n_8_57));
   NOR2_X1 i_8_0_94 (.A1(n_8_0_34), .A2(n_8_0_27), .ZN(n_8_58));
   NOR2_X1 i_8_0_95 (.A1(n_8_0_34), .A2(n_8_0_28), .ZN(n_8_59));
   NOR2_X1 i_8_0_96 (.A1(n_8_0_34), .A2(n_8_0_29), .ZN(n_8_60));
   NOR2_X1 i_8_0_97 (.A1(n_8_0_34), .A2(n_8_0_30), .ZN(n_8_61));
   NOR2_X1 i_8_0_98 (.A1(n_8_0_34), .A2(n_8_0_31), .ZN(n_8_62));
   NOR2_X1 i_8_0_99 (.A1(n_8_0_34), .A2(n_8_0_32), .ZN(n_8_63));
   NOR2_X1 i_8_0_100 (.A1(n_8_0_34), .A2(n_8_0_33), .ZN(n_8_64));
   NOR2_X1 i_8_0_103 (.A1(n_8_0_35), .A2(n_8_0_2), .ZN(n_8_66));
   NOR2_X1 i_8_0_104 (.A1(n_8_0_35), .A2(n_8_0_3), .ZN(n_8_67));
   NOR2_X1 i_8_0_105 (.A1(n_8_0_35), .A2(n_8_0_4), .ZN(n_8_68));
   NOR2_X1 i_8_0_106 (.A1(n_8_0_35), .A2(n_8_0_5), .ZN(n_8_69));
   NOR2_X1 i_8_0_107 (.A1(n_8_0_35), .A2(n_8_0_6), .ZN(n_8_70));
   NOR2_X1 i_8_0_108 (.A1(n_8_0_35), .A2(n_8_0_7), .ZN(n_8_71));
   NOR2_X1 i_8_0_109 (.A1(n_8_0_35), .A2(n_8_0_8), .ZN(n_8_72));
   NOR2_X1 i_8_0_110 (.A1(n_8_0_35), .A2(n_8_0_9), .ZN(n_8_73));
   NOR2_X1 i_8_0_111 (.A1(n_8_0_35), .A2(n_8_0_10), .ZN(n_8_74));
   NOR2_X1 i_8_0_112 (.A1(n_8_0_35), .A2(n_8_0_11), .ZN(n_8_75));
   NOR2_X1 i_8_0_113 (.A1(n_8_0_35), .A2(n_8_0_12), .ZN(n_8_76));
   NOR2_X1 i_8_0_114 (.A1(n_8_0_35), .A2(n_8_0_13), .ZN(n_8_77));
   NOR2_X1 i_8_0_115 (.A1(n_8_0_35), .A2(n_8_0_14), .ZN(n_8_78));
   NOR2_X1 i_8_0_116 (.A1(n_8_0_35), .A2(n_8_0_15), .ZN(n_8_79));
   NOR2_X1 i_8_0_117 (.A1(n_8_0_35), .A2(n_8_0_16), .ZN(n_8_80));
   NOR2_X1 i_8_0_118 (.A1(n_8_0_35), .A2(n_8_0_17), .ZN(n_8_81));
   NOR2_X1 i_8_0_119 (.A1(n_8_0_35), .A2(n_8_0_18), .ZN(n_8_82));
   NOR2_X1 i_8_0_120 (.A1(n_8_0_35), .A2(n_8_0_19), .ZN(n_8_83));
   NOR2_X1 i_8_0_121 (.A1(n_8_0_35), .A2(n_8_0_20), .ZN(n_8_84));
   NOR2_X1 i_8_0_122 (.A1(n_8_0_35), .A2(n_8_0_21), .ZN(n_8_85));
   NOR2_X1 i_8_0_123 (.A1(n_8_0_35), .A2(n_8_0_22), .ZN(n_8_86));
   NOR2_X1 i_8_0_124 (.A1(n_8_0_35), .A2(n_8_0_23), .ZN(n_8_87));
   NOR2_X1 i_8_0_125 (.A1(n_8_0_35), .A2(n_8_0_24), .ZN(n_8_88));
   NOR2_X1 i_8_0_126 (.A1(n_8_0_35), .A2(n_8_0_25), .ZN(n_8_89));
   NOR2_X1 i_8_0_127 (.A1(n_8_0_35), .A2(n_8_0_26), .ZN(n_8_90));
   NOR2_X1 i_8_0_128 (.A1(n_8_0_35), .A2(n_8_0_27), .ZN(n_8_91));
   NOR2_X1 i_8_0_129 (.A1(n_8_0_35), .A2(n_8_0_28), .ZN(n_8_92));
   NOR2_X1 i_8_0_130 (.A1(n_8_0_35), .A2(n_8_0_29), .ZN(n_8_93));
   NOR2_X1 i_8_0_131 (.A1(n_8_0_35), .A2(n_8_0_30), .ZN(n_8_94));
   NOR2_X1 i_8_0_132 (.A1(n_8_0_35), .A2(n_8_0_31), .ZN(n_8_95));
   NOR2_X1 i_8_0_133 (.A1(n_8_0_35), .A2(n_8_0_32), .ZN(n_8_96));
   NOR2_X1 i_8_0_134 (.A1(n_8_0_35), .A2(n_8_0_33), .ZN(n_8_97));
   NOR2_X1 i_8_0_139 (.A1(n_8_0_36), .A2(n_8_0_4), .ZN(n_8_101));
   NOR2_X1 i_8_0_140 (.A1(n_8_0_36), .A2(n_8_0_5), .ZN(n_8_102));
   NOR2_X1 i_8_0_141 (.A1(n_8_0_36), .A2(n_8_0_6), .ZN(n_8_103));
   NOR2_X1 i_8_0_142 (.A1(n_8_0_36), .A2(n_8_0_7), .ZN(n_8_104));
   NOR2_X1 i_8_0_143 (.A1(n_8_0_36), .A2(n_8_0_8), .ZN(n_8_105));
   NOR2_X1 i_8_0_144 (.A1(n_8_0_36), .A2(n_8_0_9), .ZN(n_8_106));
   NOR2_X1 i_8_0_145 (.A1(n_8_0_36), .A2(n_8_0_10), .ZN(n_8_107));
   NOR2_X1 i_8_0_146 (.A1(n_8_0_36), .A2(n_8_0_11), .ZN(n_8_108));
   NOR2_X1 i_8_0_147 (.A1(n_8_0_36), .A2(n_8_0_12), .ZN(n_8_109));
   NOR2_X1 i_8_0_148 (.A1(n_8_0_36), .A2(n_8_0_13), .ZN(n_8_110));
   NOR2_X1 i_8_0_149 (.A1(n_8_0_36), .A2(n_8_0_14), .ZN(n_8_111));
   NOR2_X1 i_8_0_150 (.A1(n_8_0_36), .A2(n_8_0_15), .ZN(n_8_112));
   NOR2_X1 i_8_0_151 (.A1(n_8_0_36), .A2(n_8_0_16), .ZN(n_8_113));
   NOR2_X1 i_8_0_152 (.A1(n_8_0_36), .A2(n_8_0_17), .ZN(n_8_114));
   NOR2_X1 i_8_0_153 (.A1(n_8_0_36), .A2(n_8_0_18), .ZN(n_8_115));
   NOR2_X1 i_8_0_154 (.A1(n_8_0_36), .A2(n_8_0_19), .ZN(n_8_116));
   NOR2_X1 i_8_0_155 (.A1(n_8_0_36), .A2(n_8_0_20), .ZN(n_8_117));
   NOR2_X1 i_8_0_156 (.A1(n_8_0_36), .A2(n_8_0_21), .ZN(n_8_118));
   NOR2_X1 i_8_0_157 (.A1(n_8_0_36), .A2(n_8_0_22), .ZN(n_8_119));
   NOR2_X1 i_8_0_158 (.A1(n_8_0_36), .A2(n_8_0_23), .ZN(n_8_120));
   NOR2_X1 i_8_0_159 (.A1(n_8_0_36), .A2(n_8_0_24), .ZN(n_8_121));
   NOR2_X1 i_8_0_160 (.A1(n_8_0_36), .A2(n_8_0_25), .ZN(n_8_122));
   NOR2_X1 i_8_0_161 (.A1(n_8_0_36), .A2(n_8_0_26), .ZN(n_8_123));
   NOR2_X1 i_8_0_162 (.A1(n_8_0_36), .A2(n_8_0_27), .ZN(n_8_124));
   NOR2_X1 i_8_0_163 (.A1(n_8_0_36), .A2(n_8_0_28), .ZN(n_8_125));
   NOR2_X1 i_8_0_164 (.A1(n_8_0_36), .A2(n_8_0_29), .ZN(n_8_126));
   NOR2_X1 i_8_0_165 (.A1(n_8_0_36), .A2(n_8_0_30), .ZN(n_8_127));
   NOR2_X1 i_8_0_166 (.A1(n_8_0_36), .A2(n_8_0_31), .ZN(n_8_128));
   NOR2_X1 i_8_0_167 (.A1(n_8_0_36), .A2(n_8_0_32), .ZN(n_8_129));
   NOR2_X1 i_8_0_168 (.A1(n_8_0_36), .A2(n_8_0_33), .ZN(n_8_130));
   NOR2_X1 i_8_0_171 (.A1(n_8_0_37), .A2(n_8_0_2), .ZN(n_8_132));
   NOR2_X1 i_8_0_173 (.A1(n_8_0_37), .A2(n_8_0_4), .ZN(n_8_134));
   NOR2_X1 i_8_0_174 (.A1(n_8_0_37), .A2(n_8_0_5), .ZN(n_8_135));
   NOR2_X1 i_8_0_175 (.A1(n_8_0_37), .A2(n_8_0_6), .ZN(n_8_136));
   NOR2_X1 i_8_0_176 (.A1(n_8_0_37), .A2(n_8_0_7), .ZN(n_8_137));
   NOR2_X1 i_8_0_177 (.A1(n_8_0_37), .A2(n_8_0_8), .ZN(n_8_138));
   NOR2_X1 i_8_0_178 (.A1(n_8_0_37), .A2(n_8_0_9), .ZN(n_8_139));
   NOR2_X1 i_8_0_179 (.A1(n_8_0_37), .A2(n_8_0_10), .ZN(n_8_140));
   NOR2_X1 i_8_0_180 (.A1(n_8_0_37), .A2(n_8_0_11), .ZN(n_8_141));
   NOR2_X1 i_8_0_181 (.A1(n_8_0_37), .A2(n_8_0_12), .ZN(n_8_142));
   NOR2_X1 i_8_0_182 (.A1(n_8_0_37), .A2(n_8_0_13), .ZN(n_8_143));
   NOR2_X1 i_8_0_183 (.A1(n_8_0_37), .A2(n_8_0_14), .ZN(n_8_144));
   NOR2_X1 i_8_0_184 (.A1(n_8_0_37), .A2(n_8_0_15), .ZN(n_8_145));
   NOR2_X1 i_8_0_185 (.A1(n_8_0_37), .A2(n_8_0_16), .ZN(n_8_146));
   NOR2_X1 i_8_0_186 (.A1(n_8_0_37), .A2(n_8_0_17), .ZN(n_8_147));
   NOR2_X1 i_8_0_187 (.A1(n_8_0_37), .A2(n_8_0_18), .ZN(n_8_148));
   NOR2_X1 i_8_0_188 (.A1(n_8_0_37), .A2(n_8_0_19), .ZN(n_8_149));
   NOR2_X1 i_8_0_189 (.A1(n_8_0_37), .A2(n_8_0_20), .ZN(n_8_150));
   NOR2_X1 i_8_0_190 (.A1(n_8_0_37), .A2(n_8_0_21), .ZN(n_8_151));
   NOR2_X1 i_8_0_191 (.A1(n_8_0_37), .A2(n_8_0_22), .ZN(n_8_152));
   NOR2_X1 i_8_0_192 (.A1(n_8_0_37), .A2(n_8_0_23), .ZN(n_8_153));
   NOR2_X1 i_8_0_193 (.A1(n_8_0_37), .A2(n_8_0_24), .ZN(n_8_154));
   NOR2_X1 i_8_0_194 (.A1(n_8_0_37), .A2(n_8_0_25), .ZN(n_8_155));
   NOR2_X1 i_8_0_195 (.A1(n_8_0_37), .A2(n_8_0_26), .ZN(n_8_156));
   NOR2_X1 i_8_0_196 (.A1(n_8_0_37), .A2(n_8_0_27), .ZN(n_8_157));
   NOR2_X1 i_8_0_197 (.A1(n_8_0_37), .A2(n_8_0_28), .ZN(n_8_158));
   NOR2_X1 i_8_0_198 (.A1(n_8_0_37), .A2(n_8_0_29), .ZN(n_8_159));
   NOR2_X1 i_8_0_199 (.A1(n_8_0_37), .A2(n_8_0_30), .ZN(n_8_160));
   NOR2_X1 i_8_0_200 (.A1(n_8_0_37), .A2(n_8_0_31), .ZN(n_8_161));
   NOR2_X1 i_8_0_201 (.A1(n_8_0_37), .A2(n_8_0_32), .ZN(n_8_162));
   NOR2_X1 i_8_0_202 (.A1(n_8_0_37), .A2(n_8_0_33), .ZN(n_8_163));
   NOR2_X1 i_8_0_205 (.A1(n_8_0_38), .A2(n_8_0_2), .ZN(n_8_165));
   NOR2_X1 i_8_0_206 (.A1(n_8_0_38), .A2(n_8_0_3), .ZN(n_8_166));
   NOR2_X1 i_8_0_207 (.A1(n_8_0_38), .A2(n_8_0_4), .ZN(n_8_167));
   NOR2_X1 i_8_0_208 (.A1(n_8_0_38), .A2(n_8_0_5), .ZN(n_8_168));
   NOR2_X1 i_8_0_209 (.A1(n_8_0_38), .A2(n_8_0_6), .ZN(n_8_169));
   NOR2_X1 i_8_0_210 (.A1(n_8_0_38), .A2(n_8_0_7), .ZN(n_8_170));
   NOR2_X1 i_8_0_211 (.A1(n_8_0_38), .A2(n_8_0_8), .ZN(n_8_171));
   NOR2_X1 i_8_0_212 (.A1(n_8_0_38), .A2(n_8_0_9), .ZN(n_8_172));
   NOR2_X1 i_8_0_213 (.A1(n_8_0_38), .A2(n_8_0_10), .ZN(n_8_173));
   NOR2_X1 i_8_0_214 (.A1(n_8_0_38), .A2(n_8_0_11), .ZN(n_8_174));
   NOR2_X1 i_8_0_215 (.A1(n_8_0_38), .A2(n_8_0_12), .ZN(n_8_175));
   NOR2_X1 i_8_0_216 (.A1(n_8_0_38), .A2(n_8_0_13), .ZN(n_8_176));
   NOR2_X1 i_8_0_217 (.A1(n_8_0_38), .A2(n_8_0_14), .ZN(n_8_177));
   NOR2_X1 i_8_0_218 (.A1(n_8_0_38), .A2(n_8_0_15), .ZN(n_8_178));
   NOR2_X1 i_8_0_219 (.A1(n_8_0_38), .A2(n_8_0_16), .ZN(n_8_179));
   NOR2_X1 i_8_0_220 (.A1(n_8_0_38), .A2(n_8_0_17), .ZN(n_8_180));
   NOR2_X1 i_8_0_221 (.A1(n_8_0_38), .A2(n_8_0_18), .ZN(n_8_181));
   NOR2_X1 i_8_0_222 (.A1(n_8_0_38), .A2(n_8_0_19), .ZN(n_8_182));
   NOR2_X1 i_8_0_223 (.A1(n_8_0_38), .A2(n_8_0_20), .ZN(n_8_183));
   NOR2_X1 i_8_0_224 (.A1(n_8_0_38), .A2(n_8_0_21), .ZN(n_8_184));
   NOR2_X1 i_8_0_225 (.A1(n_8_0_38), .A2(n_8_0_22), .ZN(n_8_185));
   NOR2_X1 i_8_0_226 (.A1(n_8_0_38), .A2(n_8_0_23), .ZN(n_8_186));
   NOR2_X1 i_8_0_227 (.A1(n_8_0_38), .A2(n_8_0_24), .ZN(n_8_187));
   NOR2_X1 i_8_0_228 (.A1(n_8_0_38), .A2(n_8_0_25), .ZN(n_8_188));
   NOR2_X1 i_8_0_229 (.A1(n_8_0_38), .A2(n_8_0_26), .ZN(n_8_189));
   NOR2_X1 i_8_0_230 (.A1(n_8_0_38), .A2(n_8_0_27), .ZN(n_8_190));
   NOR2_X1 i_8_0_231 (.A1(n_8_0_38), .A2(n_8_0_28), .ZN(n_8_191));
   NOR2_X1 i_8_0_232 (.A1(n_8_0_38), .A2(n_8_0_29), .ZN(n_8_192));
   NOR2_X1 i_8_0_233 (.A1(n_8_0_38), .A2(n_8_0_30), .ZN(n_8_193));
   NOR2_X1 i_8_0_234 (.A1(n_8_0_38), .A2(n_8_0_31), .ZN(n_8_194));
   NOR2_X1 i_8_0_235 (.A1(n_8_0_38), .A2(n_8_0_32), .ZN(n_8_195));
   NOR2_X1 i_8_0_236 (.A1(n_8_0_38), .A2(n_8_0_33), .ZN(n_8_196));
   NOR2_X1 i_8_0_241 (.A1(n_8_0_39), .A2(n_8_0_4), .ZN(n_8_200));
   NOR2_X1 i_8_0_242 (.A1(n_8_0_39), .A2(n_8_0_5), .ZN(n_8_201));
   NOR2_X1 i_8_0_243 (.A1(n_8_0_39), .A2(n_8_0_6), .ZN(n_8_202));
   NOR2_X1 i_8_0_244 (.A1(n_8_0_39), .A2(n_8_0_7), .ZN(n_8_203));
   NOR2_X1 i_8_0_245 (.A1(n_8_0_39), .A2(n_8_0_8), .ZN(n_8_204));
   NOR2_X1 i_8_0_246 (.A1(n_8_0_39), .A2(n_8_0_9), .ZN(n_8_205));
   NOR2_X1 i_8_0_247 (.A1(n_8_0_39), .A2(n_8_0_10), .ZN(n_8_206));
   NOR2_X1 i_8_0_248 (.A1(n_8_0_39), .A2(n_8_0_11), .ZN(n_8_207));
   NOR2_X1 i_8_0_249 (.A1(n_8_0_39), .A2(n_8_0_12), .ZN(n_8_208));
   NOR2_X1 i_8_0_250 (.A1(n_8_0_39), .A2(n_8_0_13), .ZN(n_8_209));
   NOR2_X1 i_8_0_251 (.A1(n_8_0_39), .A2(n_8_0_14), .ZN(n_8_210));
   NOR2_X1 i_8_0_252 (.A1(n_8_0_39), .A2(n_8_0_15), .ZN(n_8_211));
   NOR2_X1 i_8_0_253 (.A1(n_8_0_39), .A2(n_8_0_16), .ZN(n_8_212));
   NOR2_X1 i_8_0_254 (.A1(n_8_0_39), .A2(n_8_0_17), .ZN(n_8_213));
   NOR2_X1 i_8_0_255 (.A1(n_8_0_39), .A2(n_8_0_18), .ZN(n_8_214));
   NOR2_X1 i_8_0_256 (.A1(n_8_0_39), .A2(n_8_0_19), .ZN(n_8_215));
   NOR2_X1 i_8_0_257 (.A1(n_8_0_39), .A2(n_8_0_20), .ZN(n_8_216));
   NOR2_X1 i_8_0_258 (.A1(n_8_0_39), .A2(n_8_0_21), .ZN(n_8_217));
   NOR2_X1 i_8_0_259 (.A1(n_8_0_39), .A2(n_8_0_22), .ZN(n_8_218));
   NOR2_X1 i_8_0_260 (.A1(n_8_0_39), .A2(n_8_0_23), .ZN(n_8_219));
   NOR2_X1 i_8_0_261 (.A1(n_8_0_39), .A2(n_8_0_24), .ZN(n_8_220));
   NOR2_X1 i_8_0_262 (.A1(n_8_0_39), .A2(n_8_0_25), .ZN(n_8_221));
   NOR2_X1 i_8_0_263 (.A1(n_8_0_39), .A2(n_8_0_26), .ZN(n_8_222));
   NOR2_X1 i_8_0_264 (.A1(n_8_0_39), .A2(n_8_0_27), .ZN(n_8_223));
   NOR2_X1 i_8_0_265 (.A1(n_8_0_39), .A2(n_8_0_28), .ZN(n_8_224));
   NOR2_X1 i_8_0_266 (.A1(n_8_0_39), .A2(n_8_0_29), .ZN(n_8_225));
   NOR2_X1 i_8_0_267 (.A1(n_8_0_39), .A2(n_8_0_30), .ZN(n_8_226));
   NOR2_X1 i_8_0_268 (.A1(n_8_0_39), .A2(n_8_0_31), .ZN(n_8_227));
   NOR2_X1 i_8_0_269 (.A1(n_8_0_39), .A2(n_8_0_32), .ZN(n_8_228));
   NOR2_X1 i_8_0_270 (.A1(n_8_0_39), .A2(n_8_0_33), .ZN(n_8_229));
   NOR2_X1 i_8_0_272 (.A1(n_8_0_40), .A2(n_8_0_1), .ZN(n_8_230));
   NOR2_X1 i_8_0_277 (.A1(n_8_0_40), .A2(n_8_0_6), .ZN(n_8_235));
   NOR2_X1 i_8_0_279 (.A1(n_8_0_40), .A2(n_8_0_8), .ZN(n_8_237));
   NOR2_X1 i_8_0_281 (.A1(n_8_0_40), .A2(n_8_0_10), .ZN(n_8_239));
   NOR2_X1 i_8_0_285 (.A1(n_8_0_40), .A2(n_8_0_14), .ZN(n_8_243));
   NOR2_X1 i_8_0_286 (.A1(n_8_0_40), .A2(n_8_0_15), .ZN(n_8_244));
   NOR2_X1 i_8_0_287 (.A1(n_8_0_40), .A2(n_8_0_16), .ZN(n_8_245));
   NOR2_X1 i_8_0_288 (.A1(n_8_0_40), .A2(n_8_0_17), .ZN(n_8_246));
   NOR2_X1 i_8_0_289 (.A1(n_8_0_40), .A2(n_8_0_18), .ZN(n_8_247));
   NOR2_X1 i_8_0_290 (.A1(n_8_0_40), .A2(n_8_0_19), .ZN(n_8_248));
   NOR2_X1 i_8_0_291 (.A1(n_8_0_40), .A2(n_8_0_20), .ZN(n_8_249));
   NOR2_X1 i_8_0_292 (.A1(n_8_0_40), .A2(n_8_0_21), .ZN(n_8_250));
   NOR2_X1 i_8_0_293 (.A1(n_8_0_40), .A2(n_8_0_22), .ZN(n_8_251));
   NOR2_X1 i_8_0_294 (.A1(n_8_0_40), .A2(n_8_0_23), .ZN(n_8_252));
   NOR2_X1 i_8_0_295 (.A1(n_8_0_40), .A2(n_8_0_24), .ZN(n_8_253));
   NOR2_X1 i_8_0_296 (.A1(n_8_0_40), .A2(n_8_0_25), .ZN(n_8_254));
   NOR2_X1 i_8_0_297 (.A1(n_8_0_40), .A2(n_8_0_26), .ZN(n_8_255));
   NOR2_X1 i_8_0_298 (.A1(n_8_0_40), .A2(n_8_0_27), .ZN(n_8_256));
   NOR2_X1 i_8_0_299 (.A1(n_8_0_40), .A2(n_8_0_28), .ZN(n_8_257));
   NOR2_X1 i_8_0_300 (.A1(n_8_0_40), .A2(n_8_0_29), .ZN(n_8_258));
   NOR2_X1 i_8_0_301 (.A1(n_8_0_40), .A2(n_8_0_30), .ZN(n_8_259));
   NOR2_X1 i_8_0_302 (.A1(n_8_0_40), .A2(n_8_0_31), .ZN(n_8_260));
   NOR2_X1 i_8_0_303 (.A1(n_8_0_40), .A2(n_8_0_32), .ZN(n_8_261));
   NOR2_X1 i_8_0_304 (.A1(n_8_0_40), .A2(n_8_0_33), .ZN(n_8_262));
   INV_X1 i_8_0_305 (.A(n_102), .ZN(n_8_0_41));
   NOR2_X1 i_8_0_306 (.A1(n_8_0_41), .A2(n_8_0_1), .ZN(n_8_263));
   NOR2_X1 i_8_0_307 (.A1(n_8_0_41), .A2(n_8_0_2), .ZN(n_8_264));
   NOR2_X1 i_8_0_308 (.A1(n_8_0_41), .A2(n_8_0_3), .ZN(n_8_265));
   NOR2_X1 i_8_0_309 (.A1(n_8_0_41), .A2(n_8_0_4), .ZN(n_8_266));
   NOR2_X1 i_8_0_310 (.A1(n_8_0_41), .A2(n_8_0_5), .ZN(n_8_267));
   NOR2_X1 i_8_0_311 (.A1(n_8_0_41), .A2(n_8_0_6), .ZN(n_8_268));
   NOR2_X1 i_8_0_312 (.A1(n_8_0_41), .A2(n_8_0_7), .ZN(n_8_269));
   NOR2_X1 i_8_0_313 (.A1(n_8_0_41), .A2(n_8_0_8), .ZN(n_8_270));
   NOR2_X1 i_8_0_314 (.A1(n_8_0_41), .A2(n_8_0_9), .ZN(n_8_271));
   NOR2_X1 i_8_0_315 (.A1(n_8_0_41), .A2(n_8_0_10), .ZN(n_8_272));
   NOR2_X1 i_8_0_316 (.A1(n_8_0_41), .A2(n_8_0_11), .ZN(n_8_273));
   NOR2_X1 i_8_0_317 (.A1(n_8_0_41), .A2(n_8_0_12), .ZN(n_8_274));
   NOR2_X1 i_8_0_318 (.A1(n_8_0_41), .A2(n_8_0_13), .ZN(n_8_275));
   NOR2_X1 i_8_0_319 (.A1(n_8_0_41), .A2(n_8_0_14), .ZN(n_8_276));
   NOR2_X1 i_8_0_320 (.A1(n_8_0_41), .A2(n_8_0_15), .ZN(n_8_277));
   NOR2_X1 i_8_0_321 (.A1(n_8_0_41), .A2(n_8_0_16), .ZN(n_8_278));
   NOR2_X1 i_8_0_322 (.A1(n_8_0_41), .A2(n_8_0_17), .ZN(n_8_279));
   NOR2_X1 i_8_0_323 (.A1(n_8_0_41), .A2(n_8_0_18), .ZN(n_8_280));
   NOR2_X1 i_8_0_324 (.A1(n_8_0_41), .A2(n_8_0_19), .ZN(n_8_281));
   NOR2_X1 i_8_0_325 (.A1(n_8_0_41), .A2(n_8_0_20), .ZN(n_8_282));
   NOR2_X1 i_8_0_326 (.A1(n_8_0_41), .A2(n_8_0_21), .ZN(n_8_283));
   NOR2_X1 i_8_0_327 (.A1(n_8_0_41), .A2(n_8_0_22), .ZN(n_8_284));
   NOR2_X1 i_8_0_328 (.A1(n_8_0_41), .A2(n_8_0_23), .ZN(n_8_285));
   NOR2_X1 i_8_0_329 (.A1(n_8_0_41), .A2(n_8_0_24), .ZN(n_8_286));
   NOR2_X1 i_8_0_330 (.A1(n_8_0_41), .A2(n_8_0_25), .ZN(n_8_287));
   NOR2_X1 i_8_0_331 (.A1(n_8_0_41), .A2(n_8_0_26), .ZN(n_8_288));
   NOR2_X1 i_8_0_332 (.A1(n_8_0_41), .A2(n_8_0_27), .ZN(n_8_289));
   NOR2_X1 i_8_0_333 (.A1(n_8_0_41), .A2(n_8_0_28), .ZN(n_8_290));
   NOR2_X1 i_8_0_334 (.A1(n_8_0_41), .A2(n_8_0_29), .ZN(n_8_291));
   NOR2_X1 i_8_0_335 (.A1(n_8_0_41), .A2(n_8_0_30), .ZN(n_8_292));
   NOR2_X1 i_8_0_336 (.A1(n_8_0_41), .A2(n_8_0_31), .ZN(n_8_293));
   NOR2_X1 i_8_0_337 (.A1(n_8_0_41), .A2(n_8_0_32), .ZN(n_8_294));
   NOR2_X1 i_8_0_338 (.A1(n_8_0_41), .A2(n_8_0_33), .ZN(n_8_295));
   INV_X1 i_8_0_339 (.A(n_78), .ZN(n_8_0_42));
   NOR2_X1 i_8_0_340 (.A1(n_8_0_42), .A2(n_8_0_1), .ZN(n_8_296));
   NOR2_X1 i_8_0_341 (.A1(n_8_0_42), .A2(n_8_0_2), .ZN(n_8_297));
   NOR2_X1 i_8_0_342 (.A1(n_8_0_42), .A2(n_8_0_3), .ZN(n_8_298));
   NOR2_X1 i_8_0_343 (.A1(n_8_0_42), .A2(n_8_0_4), .ZN(n_8_299));
   NOR2_X1 i_8_0_344 (.A1(n_8_0_42), .A2(n_8_0_5), .ZN(n_8_300));
   NOR2_X1 i_8_0_345 (.A1(n_8_0_42), .A2(n_8_0_6), .ZN(n_8_301));
   NOR2_X1 i_8_0_346 (.A1(n_8_0_42), .A2(n_8_0_7), .ZN(n_8_302));
   NOR2_X1 i_8_0_347 (.A1(n_8_0_42), .A2(n_8_0_8), .ZN(n_8_303));
   NOR2_X1 i_8_0_348 (.A1(n_8_0_42), .A2(n_8_0_9), .ZN(n_8_304));
   NOR2_X1 i_8_0_349 (.A1(n_8_0_42), .A2(n_8_0_10), .ZN(n_8_305));
   NOR2_X1 i_8_0_350 (.A1(n_8_0_42), .A2(n_8_0_11), .ZN(n_8_306));
   NOR2_X1 i_8_0_351 (.A1(n_8_0_42), .A2(n_8_0_12), .ZN(n_8_307));
   NOR2_X1 i_8_0_352 (.A1(n_8_0_42), .A2(n_8_0_13), .ZN(n_8_308));
   NOR2_X1 i_8_0_353 (.A1(n_8_0_42), .A2(n_8_0_14), .ZN(n_8_309));
   NOR2_X1 i_8_0_354 (.A1(n_8_0_42), .A2(n_8_0_15), .ZN(n_8_310));
   NOR2_X1 i_8_0_355 (.A1(n_8_0_42), .A2(n_8_0_16), .ZN(n_8_311));
   NOR2_X1 i_8_0_356 (.A1(n_8_0_42), .A2(n_8_0_17), .ZN(n_8_312));
   NOR2_X1 i_8_0_357 (.A1(n_8_0_42), .A2(n_8_0_18), .ZN(n_8_313));
   NOR2_X1 i_8_0_358 (.A1(n_8_0_42), .A2(n_8_0_19), .ZN(n_8_314));
   NOR2_X1 i_8_0_359 (.A1(n_8_0_42), .A2(n_8_0_20), .ZN(n_8_315));
   NOR2_X1 i_8_0_360 (.A1(n_8_0_42), .A2(n_8_0_21), .ZN(n_8_316));
   NOR2_X1 i_8_0_361 (.A1(n_8_0_42), .A2(n_8_0_22), .ZN(n_8_317));
   NOR2_X1 i_8_0_362 (.A1(n_8_0_42), .A2(n_8_0_23), .ZN(n_8_318));
   NOR2_X1 i_8_0_363 (.A1(n_8_0_42), .A2(n_8_0_24), .ZN(n_8_319));
   NOR2_X1 i_8_0_364 (.A1(n_8_0_42), .A2(n_8_0_25), .ZN(n_8_320));
   NOR2_X1 i_8_0_365 (.A1(n_8_0_42), .A2(n_8_0_26), .ZN(n_8_321));
   NOR2_X1 i_8_0_366 (.A1(n_8_0_42), .A2(n_8_0_27), .ZN(n_8_322));
   NOR2_X1 i_8_0_367 (.A1(n_8_0_42), .A2(n_8_0_28), .ZN(n_8_323));
   NOR2_X1 i_8_0_368 (.A1(n_8_0_42), .A2(n_8_0_29), .ZN(n_8_324));
   NOR2_X1 i_8_0_369 (.A1(n_8_0_42), .A2(n_8_0_30), .ZN(n_8_325));
   NOR2_X1 i_8_0_370 (.A1(n_8_0_42), .A2(n_8_0_31), .ZN(n_8_326));
   NOR2_X1 i_8_0_371 (.A1(n_8_0_42), .A2(n_8_0_32), .ZN(n_8_327));
   NOR2_X1 i_8_0_372 (.A1(n_8_0_42), .A2(n_8_0_33), .ZN(n_8_328));
   INV_X1 i_8_0_373 (.A(n_101), .ZN(n_8_0_43));
   NOR2_X1 i_8_0_374 (.A1(n_8_0_43), .A2(n_8_0_1), .ZN(n_8_329));
   NOR2_X1 i_8_0_375 (.A1(n_8_0_43), .A2(n_8_0_2), .ZN(n_8_330));
   NOR2_X1 i_8_0_376 (.A1(n_8_0_43), .A2(n_8_0_3), .ZN(n_8_331));
   NOR2_X1 i_8_0_377 (.A1(n_8_0_43), .A2(n_8_0_4), .ZN(n_8_332));
   NOR2_X1 i_8_0_378 (.A1(n_8_0_43), .A2(n_8_0_5), .ZN(n_8_333));
   NOR2_X1 i_8_0_379 (.A1(n_8_0_43), .A2(n_8_0_6), .ZN(n_8_334));
   NOR2_X1 i_8_0_380 (.A1(n_8_0_43), .A2(n_8_0_7), .ZN(n_8_335));
   NOR2_X1 i_8_0_381 (.A1(n_8_0_43), .A2(n_8_0_8), .ZN(n_8_336));
   NOR2_X1 i_8_0_382 (.A1(n_8_0_43), .A2(n_8_0_9), .ZN(n_8_337));
   NOR2_X1 i_8_0_383 (.A1(n_8_0_43), .A2(n_8_0_10), .ZN(n_8_338));
   NOR2_X1 i_8_0_384 (.A1(n_8_0_43), .A2(n_8_0_11), .ZN(n_8_339));
   NOR2_X1 i_8_0_385 (.A1(n_8_0_43), .A2(n_8_0_12), .ZN(n_8_340));
   NOR2_X1 i_8_0_386 (.A1(n_8_0_43), .A2(n_8_0_13), .ZN(n_8_341));
   NOR2_X1 i_8_0_387 (.A1(n_8_0_43), .A2(n_8_0_14), .ZN(n_8_342));
   NOR2_X1 i_8_0_388 (.A1(n_8_0_43), .A2(n_8_0_15), .ZN(n_8_343));
   NOR2_X1 i_8_0_389 (.A1(n_8_0_43), .A2(n_8_0_16), .ZN(n_8_344));
   NOR2_X1 i_8_0_390 (.A1(n_8_0_43), .A2(n_8_0_17), .ZN(n_8_345));
   NOR2_X1 i_8_0_391 (.A1(n_8_0_43), .A2(n_8_0_18), .ZN(n_8_346));
   NOR2_X1 i_8_0_392 (.A1(n_8_0_43), .A2(n_8_0_19), .ZN(n_8_347));
   NOR2_X1 i_8_0_393 (.A1(n_8_0_43), .A2(n_8_0_20), .ZN(n_8_348));
   NOR2_X1 i_8_0_394 (.A1(n_8_0_43), .A2(n_8_0_21), .ZN(n_8_349));
   NOR2_X1 i_8_0_395 (.A1(n_8_0_43), .A2(n_8_0_22), .ZN(n_8_350));
   NOR2_X1 i_8_0_396 (.A1(n_8_0_43), .A2(n_8_0_23), .ZN(n_8_351));
   NOR2_X1 i_8_0_397 (.A1(n_8_0_43), .A2(n_8_0_24), .ZN(n_8_352));
   NOR2_X1 i_8_0_398 (.A1(n_8_0_43), .A2(n_8_0_25), .ZN(n_8_353));
   NOR2_X1 i_8_0_399 (.A1(n_8_0_43), .A2(n_8_0_26), .ZN(n_8_354));
   NOR2_X1 i_8_0_400 (.A1(n_8_0_43), .A2(n_8_0_27), .ZN(n_8_355));
   NOR2_X1 i_8_0_401 (.A1(n_8_0_43), .A2(n_8_0_28), .ZN(n_8_356));
   NOR2_X1 i_8_0_402 (.A1(n_8_0_43), .A2(n_8_0_29), .ZN(n_8_357));
   NOR2_X1 i_8_0_403 (.A1(n_8_0_43), .A2(n_8_0_30), .ZN(n_8_358));
   NOR2_X1 i_8_0_404 (.A1(n_8_0_43), .A2(n_8_0_31), .ZN(n_8_359));
   NOR2_X1 i_8_0_405 (.A1(n_8_0_43), .A2(n_8_0_32), .ZN(n_8_360));
   NOR2_X1 i_8_0_406 (.A1(n_8_0_43), .A2(n_8_0_33), .ZN(n_8_361));
   INV_X1 i_8_0_407 (.A(n_100), .ZN(n_8_0_44));
   NOR2_X1 i_8_0_408 (.A1(n_8_0_44), .A2(n_8_0_1), .ZN(n_8_362));
   NOR2_X1 i_8_0_409 (.A1(n_8_0_44), .A2(n_8_0_2), .ZN(n_8_363));
   NOR2_X1 i_8_0_410 (.A1(n_8_0_44), .A2(n_8_0_3), .ZN(n_8_364));
   NOR2_X1 i_8_0_411 (.A1(n_8_0_44), .A2(n_8_0_4), .ZN(n_8_365));
   NOR2_X1 i_8_0_412 (.A1(n_8_0_44), .A2(n_8_0_5), .ZN(n_8_366));
   NOR2_X1 i_8_0_413 (.A1(n_8_0_44), .A2(n_8_0_6), .ZN(n_8_367));
   NOR2_X1 i_8_0_414 (.A1(n_8_0_44), .A2(n_8_0_7), .ZN(n_8_368));
   NOR2_X1 i_8_0_415 (.A1(n_8_0_44), .A2(n_8_0_8), .ZN(n_8_369));
   NOR2_X1 i_8_0_416 (.A1(n_8_0_44), .A2(n_8_0_9), .ZN(n_8_370));
   NOR2_X1 i_8_0_417 (.A1(n_8_0_44), .A2(n_8_0_10), .ZN(n_8_371));
   NOR2_X1 i_8_0_418 (.A1(n_8_0_44), .A2(n_8_0_11), .ZN(n_8_372));
   NOR2_X1 i_8_0_419 (.A1(n_8_0_44), .A2(n_8_0_12), .ZN(n_8_373));
   NOR2_X1 i_8_0_420 (.A1(n_8_0_44), .A2(n_8_0_13), .ZN(n_8_374));
   NOR2_X1 i_8_0_421 (.A1(n_8_0_44), .A2(n_8_0_14), .ZN(n_8_375));
   NOR2_X1 i_8_0_422 (.A1(n_8_0_44), .A2(n_8_0_15), .ZN(n_8_376));
   NOR2_X1 i_8_0_423 (.A1(n_8_0_44), .A2(n_8_0_16), .ZN(n_8_377));
   NOR2_X1 i_8_0_424 (.A1(n_8_0_44), .A2(n_8_0_17), .ZN(n_8_378));
   NOR2_X1 i_8_0_425 (.A1(n_8_0_44), .A2(n_8_0_18), .ZN(n_8_379));
   NOR2_X1 i_8_0_426 (.A1(n_8_0_44), .A2(n_8_0_19), .ZN(n_8_380));
   NOR2_X1 i_8_0_427 (.A1(n_8_0_44), .A2(n_8_0_20), .ZN(n_8_381));
   NOR2_X1 i_8_0_428 (.A1(n_8_0_44), .A2(n_8_0_21), .ZN(n_8_382));
   NOR2_X1 i_8_0_429 (.A1(n_8_0_44), .A2(n_8_0_22), .ZN(n_8_383));
   NOR2_X1 i_8_0_430 (.A1(n_8_0_44), .A2(n_8_0_23), .ZN(n_8_384));
   NOR2_X1 i_8_0_431 (.A1(n_8_0_44), .A2(n_8_0_24), .ZN(n_8_385));
   NOR2_X1 i_8_0_432 (.A1(n_8_0_44), .A2(n_8_0_25), .ZN(n_8_386));
   NOR2_X1 i_8_0_433 (.A1(n_8_0_44), .A2(n_8_0_26), .ZN(n_8_387));
   NOR2_X1 i_8_0_434 (.A1(n_8_0_44), .A2(n_8_0_27), .ZN(n_8_388));
   NOR2_X1 i_8_0_435 (.A1(n_8_0_44), .A2(n_8_0_28), .ZN(n_8_389));
   NOR2_X1 i_8_0_436 (.A1(n_8_0_44), .A2(n_8_0_29), .ZN(n_8_390));
   NOR2_X1 i_8_0_437 (.A1(n_8_0_44), .A2(n_8_0_30), .ZN(n_8_391));
   NOR2_X1 i_8_0_438 (.A1(n_8_0_44), .A2(n_8_0_31), .ZN(n_8_392));
   NOR2_X1 i_8_0_439 (.A1(n_8_0_44), .A2(n_8_0_32), .ZN(n_8_393));
   NOR2_X1 i_8_0_440 (.A1(n_8_0_44), .A2(n_8_0_33), .ZN(n_8_394));
   INV_X1 i_8_0_441 (.A(n_99), .ZN(n_8_0_45));
   NOR2_X1 i_8_0_442 (.A1(n_8_0_45), .A2(n_8_0_1), .ZN(n_8_1026));
   NOR2_X1 i_8_0_443 (.A1(n_8_0_45), .A2(n_8_0_2), .ZN(n_8_1027));
   NOR2_X1 i_8_0_444 (.A1(n_8_0_45), .A2(n_8_0_3), .ZN(n_8_1028));
   NOR2_X1 i_8_0_445 (.A1(n_8_0_45), .A2(n_8_0_4), .ZN(n_8_1029));
   NOR2_X1 i_8_0_446 (.A1(n_8_0_45), .A2(n_8_0_5), .ZN(n_8_1030));
   NOR2_X1 i_8_0_447 (.A1(n_8_0_45), .A2(n_8_0_6), .ZN(n_8_1031));
   NOR2_X1 i_8_0_448 (.A1(n_8_0_45), .A2(n_8_0_7), .ZN(n_8_1032));
   NOR2_X1 i_8_0_449 (.A1(n_8_0_45), .A2(n_8_0_8), .ZN(n_8_1033));
   NOR2_X1 i_8_0_450 (.A1(n_8_0_45), .A2(n_8_0_9), .ZN(n_8_1034));
   NOR2_X1 i_8_0_451 (.A1(n_8_0_45), .A2(n_8_0_10), .ZN(n_8_1035));
   NOR2_X1 i_8_0_452 (.A1(n_8_0_45), .A2(n_8_0_11), .ZN(n_8_1036));
   NOR2_X1 i_8_0_453 (.A1(n_8_0_45), .A2(n_8_0_12), .ZN(n_8_1037));
   NOR2_X1 i_8_0_454 (.A1(n_8_0_45), .A2(n_8_0_13), .ZN(n_8_1038));
   NOR2_X1 i_8_0_455 (.A1(n_8_0_45), .A2(n_8_0_14), .ZN(n_8_1039));
   NOR2_X1 i_8_0_456 (.A1(n_8_0_45), .A2(n_8_0_15), .ZN(n_8_1040));
   NOR2_X1 i_8_0_457 (.A1(n_8_0_45), .A2(n_8_0_16), .ZN(n_8_1041));
   NOR2_X1 i_8_0_458 (.A1(n_8_0_45), .A2(n_8_0_17), .ZN(n_8_1042));
   NOR2_X1 i_8_0_459 (.A1(n_8_0_45), .A2(n_8_0_18), .ZN(n_8_1043));
   NOR2_X1 i_8_0_460 (.A1(n_8_0_45), .A2(n_8_0_19), .ZN(n_8_1044));
   NOR2_X1 i_8_0_461 (.A1(n_8_0_45), .A2(n_8_0_20), .ZN(n_8_1045));
   NOR2_X1 i_8_0_462 (.A1(n_8_0_45), .A2(n_8_0_21), .ZN(n_8_1046));
   NOR2_X1 i_8_0_463 (.A1(n_8_0_45), .A2(n_8_0_22), .ZN(n_8_1047));
   NOR2_X1 i_8_0_464 (.A1(n_8_0_45), .A2(n_8_0_23), .ZN(n_8_1048));
   NOR2_X1 i_8_0_465 (.A1(n_8_0_45), .A2(n_8_0_24), .ZN(n_8_1049));
   NOR2_X1 i_8_0_466 (.A1(n_8_0_45), .A2(n_8_0_25), .ZN(n_8_1050));
   NOR2_X1 i_8_0_467 (.A1(n_8_0_45), .A2(n_8_0_26), .ZN(n_8_1051));
   NOR2_X1 i_8_0_468 (.A1(n_8_0_45), .A2(n_8_0_27), .ZN(n_8_1052));
   NOR2_X1 i_8_0_469 (.A1(n_8_0_45), .A2(n_8_0_28), .ZN(n_8_1053));
   NOR2_X1 i_8_0_470 (.A1(n_8_0_45), .A2(n_8_0_29), .ZN(n_8_1054));
   NOR2_X1 i_8_0_471 (.A1(n_8_0_45), .A2(n_8_0_30), .ZN(n_8_395));
   NOR2_X1 i_8_0_472 (.A1(n_8_0_45), .A2(n_8_0_31), .ZN(n_8_396));
   NOR2_X1 i_8_0_473 (.A1(n_8_0_45), .A2(n_8_0_32), .ZN(n_8_397));
   NOR2_X1 i_8_0_474 (.A1(n_8_0_45), .A2(n_8_0_33), .ZN(n_8_398));
   INV_X1 i_8_0_475 (.A(n_98), .ZN(n_8_0_46));
   NOR2_X1 i_8_0_476 (.A1(n_8_0_46), .A2(n_8_0_1), .ZN(n_8_981));
   NOR2_X1 i_8_0_477 (.A1(n_8_0_46), .A2(n_8_0_2), .ZN(n_8_982));
   NOR2_X1 i_8_0_478 (.A1(n_8_0_46), .A2(n_8_0_3), .ZN(n_8_983));
   NOR2_X1 i_8_0_479 (.A1(n_8_0_46), .A2(n_8_0_4), .ZN(n_8_984));
   NOR2_X1 i_8_0_480 (.A1(n_8_0_46), .A2(n_8_0_5), .ZN(n_8_985));
   NOR2_X1 i_8_0_481 (.A1(n_8_0_46), .A2(n_8_0_6), .ZN(n_8_986));
   NOR2_X1 i_8_0_482 (.A1(n_8_0_46), .A2(n_8_0_7), .ZN(n_8_987));
   NOR2_X1 i_8_0_483 (.A1(n_8_0_46), .A2(n_8_0_8), .ZN(n_8_988));
   NOR2_X1 i_8_0_484 (.A1(n_8_0_46), .A2(n_8_0_9), .ZN(n_8_989));
   NOR2_X1 i_8_0_485 (.A1(n_8_0_46), .A2(n_8_0_10), .ZN(n_8_990));
   NOR2_X1 i_8_0_486 (.A1(n_8_0_46), .A2(n_8_0_11), .ZN(n_8_991));
   NOR2_X1 i_8_0_487 (.A1(n_8_0_46), .A2(n_8_0_12), .ZN(n_8_992));
   NOR2_X1 i_8_0_488 (.A1(n_8_0_46), .A2(n_8_0_13), .ZN(n_8_993));
   NOR2_X1 i_8_0_489 (.A1(n_8_0_46), .A2(n_8_0_14), .ZN(n_8_994));
   NOR2_X1 i_8_0_490 (.A1(n_8_0_46), .A2(n_8_0_15), .ZN(n_8_995));
   NOR2_X1 i_8_0_491 (.A1(n_8_0_46), .A2(n_8_0_16), .ZN(n_8_996));
   NOR2_X1 i_8_0_492 (.A1(n_8_0_46), .A2(n_8_0_17), .ZN(n_8_997));
   NOR2_X1 i_8_0_493 (.A1(n_8_0_46), .A2(n_8_0_18), .ZN(n_8_998));
   NOR2_X1 i_8_0_494 (.A1(n_8_0_46), .A2(n_8_0_19), .ZN(n_8_999));
   NOR2_X1 i_8_0_495 (.A1(n_8_0_46), .A2(n_8_0_20), .ZN(n_8_1000));
   NOR2_X1 i_8_0_496 (.A1(n_8_0_46), .A2(n_8_0_21), .ZN(n_8_1001));
   NOR2_X1 i_8_0_497 (.A1(n_8_0_46), .A2(n_8_0_22), .ZN(n_8_1002));
   NOR2_X1 i_8_0_498 (.A1(n_8_0_46), .A2(n_8_0_23), .ZN(n_8_1003));
   NOR2_X1 i_8_0_499 (.A1(n_8_0_46), .A2(n_8_0_24), .ZN(n_8_1004));
   NOR2_X1 i_8_0_500 (.A1(n_8_0_46), .A2(n_8_0_25), .ZN(n_8_1005));
   NOR2_X1 i_8_0_501 (.A1(n_8_0_46), .A2(n_8_0_26), .ZN(n_8_1006));
   NOR2_X1 i_8_0_502 (.A1(n_8_0_46), .A2(n_8_0_27), .ZN(n_8_1007));
   NOR2_X1 i_8_0_503 (.A1(n_8_0_46), .A2(n_8_0_28), .ZN(n_8_1008));
   NOR2_X1 i_8_0_504 (.A1(n_8_0_46), .A2(n_8_0_29), .ZN(n_8_1009));
   NOR2_X1 i_8_0_505 (.A1(n_8_0_46), .A2(n_8_0_30), .ZN(n_8_1010));
   NOR2_X1 i_8_0_506 (.A1(n_8_0_46), .A2(n_8_0_31), .ZN(n_8_1011));
   NOR2_X1 i_8_0_507 (.A1(n_8_0_46), .A2(n_8_0_32), .ZN(n_8_1012));
   NOR2_X1 i_8_0_508 (.A1(n_8_0_46), .A2(n_8_0_33), .ZN(n_8_1024));
   INV_X1 i_8_0_509 (.A(n_97), .ZN(n_8_0_47));
   NOR2_X1 i_8_0_510 (.A1(n_8_0_47), .A2(n_8_0_1), .ZN(n_8_935));
   NOR2_X1 i_8_0_511 (.A1(n_8_0_47), .A2(n_8_0_2), .ZN(n_8_936));
   NOR2_X1 i_8_0_512 (.A1(n_8_0_47), .A2(n_8_0_3), .ZN(n_8_937));
   NOR2_X1 i_8_0_513 (.A1(n_8_0_47), .A2(n_8_0_4), .ZN(n_8_938));
   NOR2_X1 i_8_0_514 (.A1(n_8_0_47), .A2(n_8_0_5), .ZN(n_8_939));
   NOR2_X1 i_8_0_515 (.A1(n_8_0_47), .A2(n_8_0_6), .ZN(n_8_940));
   NOR2_X1 i_8_0_516 (.A1(n_8_0_47), .A2(n_8_0_7), .ZN(n_8_941));
   NOR2_X1 i_8_0_517 (.A1(n_8_0_47), .A2(n_8_0_8), .ZN(n_8_942));
   NOR2_X1 i_8_0_518 (.A1(n_8_0_47), .A2(n_8_0_9), .ZN(n_8_943));
   NOR2_X1 i_8_0_519 (.A1(n_8_0_47), .A2(n_8_0_10), .ZN(n_8_944));
   NOR2_X1 i_8_0_520 (.A1(n_8_0_47), .A2(n_8_0_11), .ZN(n_8_945));
   NOR2_X1 i_8_0_521 (.A1(n_8_0_47), .A2(n_8_0_12), .ZN(n_8_946));
   NOR2_X1 i_8_0_522 (.A1(n_8_0_47), .A2(n_8_0_13), .ZN(n_8_947));
   NOR2_X1 i_8_0_523 (.A1(n_8_0_47), .A2(n_8_0_14), .ZN(n_8_948));
   NOR2_X1 i_8_0_524 (.A1(n_8_0_47), .A2(n_8_0_15), .ZN(n_8_949));
   NOR2_X1 i_8_0_525 (.A1(n_8_0_47), .A2(n_8_0_16), .ZN(n_8_950));
   NOR2_X1 i_8_0_526 (.A1(n_8_0_47), .A2(n_8_0_17), .ZN(n_8_951));
   NOR2_X1 i_8_0_527 (.A1(n_8_0_47), .A2(n_8_0_18), .ZN(n_8_952));
   NOR2_X1 i_8_0_528 (.A1(n_8_0_47), .A2(n_8_0_19), .ZN(n_8_953));
   NOR2_X1 i_8_0_529 (.A1(n_8_0_47), .A2(n_8_0_20), .ZN(n_8_954));
   NOR2_X1 i_8_0_530 (.A1(n_8_0_47), .A2(n_8_0_21), .ZN(n_8_955));
   NOR2_X1 i_8_0_531 (.A1(n_8_0_47), .A2(n_8_0_22), .ZN(n_8_956));
   NOR2_X1 i_8_0_532 (.A1(n_8_0_47), .A2(n_8_0_23), .ZN(n_8_957));
   NOR2_X1 i_8_0_533 (.A1(n_8_0_47), .A2(n_8_0_24), .ZN(n_8_958));
   NOR2_X1 i_8_0_534 (.A1(n_8_0_47), .A2(n_8_0_25), .ZN(n_8_959));
   NOR2_X1 i_8_0_535 (.A1(n_8_0_47), .A2(n_8_0_26), .ZN(n_8_960));
   NOR2_X1 i_8_0_536 (.A1(n_8_0_47), .A2(n_8_0_27), .ZN(n_8_961));
   NOR2_X1 i_8_0_537 (.A1(n_8_0_47), .A2(n_8_0_28), .ZN(n_8_962));
   NOR2_X1 i_8_0_538 (.A1(n_8_0_47), .A2(n_8_0_29), .ZN(n_8_963));
   NOR2_X1 i_8_0_539 (.A1(n_8_0_47), .A2(n_8_0_30), .ZN(n_8_964));
   NOR2_X1 i_8_0_540 (.A1(n_8_0_47), .A2(n_8_0_31), .ZN(n_8_965));
   NOR2_X1 i_8_0_541 (.A1(n_8_0_47), .A2(n_8_0_32), .ZN(n_8_966));
   NOR2_X1 i_8_0_542 (.A1(n_8_0_47), .A2(n_8_0_33), .ZN(n_8_979));
   INV_X1 i_8_0_543 (.A(n_96), .ZN(n_8_0_48));
   NOR2_X1 i_8_0_544 (.A1(n_8_0_48), .A2(n_8_0_1), .ZN(n_8_888));
   NOR2_X1 i_8_0_545 (.A1(n_8_0_48), .A2(n_8_0_2), .ZN(n_8_889));
   NOR2_X1 i_8_0_546 (.A1(n_8_0_48), .A2(n_8_0_3), .ZN(n_8_890));
   NOR2_X1 i_8_0_547 (.A1(n_8_0_48), .A2(n_8_0_4), .ZN(n_8_891));
   NOR2_X1 i_8_0_548 (.A1(n_8_0_48), .A2(n_8_0_5), .ZN(n_8_892));
   NOR2_X1 i_8_0_549 (.A1(n_8_0_48), .A2(n_8_0_6), .ZN(n_8_893));
   NOR2_X1 i_8_0_550 (.A1(n_8_0_48), .A2(n_8_0_7), .ZN(n_8_894));
   NOR2_X1 i_8_0_551 (.A1(n_8_0_48), .A2(n_8_0_8), .ZN(n_8_895));
   NOR2_X1 i_8_0_552 (.A1(n_8_0_48), .A2(n_8_0_9), .ZN(n_8_896));
   NOR2_X1 i_8_0_553 (.A1(n_8_0_48), .A2(n_8_0_10), .ZN(n_8_897));
   NOR2_X1 i_8_0_554 (.A1(n_8_0_48), .A2(n_8_0_11), .ZN(n_8_898));
   NOR2_X1 i_8_0_555 (.A1(n_8_0_48), .A2(n_8_0_12), .ZN(n_8_899));
   NOR2_X1 i_8_0_556 (.A1(n_8_0_48), .A2(n_8_0_13), .ZN(n_8_900));
   NOR2_X1 i_8_0_557 (.A1(n_8_0_48), .A2(n_8_0_14), .ZN(n_8_901));
   NOR2_X1 i_8_0_558 (.A1(n_8_0_48), .A2(n_8_0_15), .ZN(n_8_902));
   NOR2_X1 i_8_0_559 (.A1(n_8_0_48), .A2(n_8_0_16), .ZN(n_8_903));
   NOR2_X1 i_8_0_560 (.A1(n_8_0_48), .A2(n_8_0_17), .ZN(n_8_904));
   NOR2_X1 i_8_0_561 (.A1(n_8_0_48), .A2(n_8_0_18), .ZN(n_8_905));
   NOR2_X1 i_8_0_562 (.A1(n_8_0_48), .A2(n_8_0_19), .ZN(n_8_906));
   NOR2_X1 i_8_0_563 (.A1(n_8_0_48), .A2(n_8_0_20), .ZN(n_8_907));
   NOR2_X1 i_8_0_564 (.A1(n_8_0_48), .A2(n_8_0_21), .ZN(n_8_908));
   NOR2_X1 i_8_0_565 (.A1(n_8_0_48), .A2(n_8_0_22), .ZN(n_8_909));
   NOR2_X1 i_8_0_566 (.A1(n_8_0_48), .A2(n_8_0_23), .ZN(n_8_910));
   NOR2_X1 i_8_0_567 (.A1(n_8_0_48), .A2(n_8_0_24), .ZN(n_8_911));
   NOR2_X1 i_8_0_568 (.A1(n_8_0_48), .A2(n_8_0_25), .ZN(n_8_912));
   NOR2_X1 i_8_0_569 (.A1(n_8_0_48), .A2(n_8_0_26), .ZN(n_8_913));
   NOR2_X1 i_8_0_570 (.A1(n_8_0_48), .A2(n_8_0_27), .ZN(n_8_914));
   NOR2_X1 i_8_0_571 (.A1(n_8_0_48), .A2(n_8_0_28), .ZN(n_8_915));
   NOR2_X1 i_8_0_572 (.A1(n_8_0_48), .A2(n_8_0_29), .ZN(n_8_916));
   NOR2_X1 i_8_0_573 (.A1(n_8_0_48), .A2(n_8_0_30), .ZN(n_8_917));
   NOR2_X1 i_8_0_574 (.A1(n_8_0_48), .A2(n_8_0_31), .ZN(n_8_918));
   NOR2_X1 i_8_0_575 (.A1(n_8_0_48), .A2(n_8_0_32), .ZN(n_8_919));
   NOR2_X1 i_8_0_576 (.A1(n_8_0_48), .A2(n_8_0_33), .ZN(n_8_933));
   INV_X1 i_8_0_577 (.A(n_95), .ZN(n_8_0_49));
   NOR2_X1 i_8_0_578 (.A1(n_8_0_49), .A2(n_8_0_1), .ZN(n_8_840));
   NOR2_X1 i_8_0_579 (.A1(n_8_0_49), .A2(n_8_0_2), .ZN(n_8_841));
   NOR2_X1 i_8_0_580 (.A1(n_8_0_49), .A2(n_8_0_3), .ZN(n_8_842));
   NOR2_X1 i_8_0_581 (.A1(n_8_0_49), .A2(n_8_0_4), .ZN(n_8_843));
   NOR2_X1 i_8_0_582 (.A1(n_8_0_49), .A2(n_8_0_5), .ZN(n_8_844));
   NOR2_X1 i_8_0_583 (.A1(n_8_0_49), .A2(n_8_0_6), .ZN(n_8_845));
   NOR2_X1 i_8_0_584 (.A1(n_8_0_49), .A2(n_8_0_7), .ZN(n_8_846));
   NOR2_X1 i_8_0_585 (.A1(n_8_0_49), .A2(n_8_0_8), .ZN(n_8_847));
   NOR2_X1 i_8_0_586 (.A1(n_8_0_49), .A2(n_8_0_9), .ZN(n_8_848));
   NOR2_X1 i_8_0_587 (.A1(n_8_0_49), .A2(n_8_0_10), .ZN(n_8_849));
   NOR2_X1 i_8_0_588 (.A1(n_8_0_49), .A2(n_8_0_11), .ZN(n_8_850));
   NOR2_X1 i_8_0_589 (.A1(n_8_0_49), .A2(n_8_0_12), .ZN(n_8_851));
   NOR2_X1 i_8_0_590 (.A1(n_8_0_49), .A2(n_8_0_13), .ZN(n_8_852));
   NOR2_X1 i_8_0_591 (.A1(n_8_0_49), .A2(n_8_0_14), .ZN(n_8_853));
   NOR2_X1 i_8_0_592 (.A1(n_8_0_49), .A2(n_8_0_15), .ZN(n_8_854));
   NOR2_X1 i_8_0_593 (.A1(n_8_0_49), .A2(n_8_0_16), .ZN(n_8_855));
   NOR2_X1 i_8_0_594 (.A1(n_8_0_49), .A2(n_8_0_17), .ZN(n_8_856));
   NOR2_X1 i_8_0_595 (.A1(n_8_0_49), .A2(n_8_0_18), .ZN(n_8_857));
   NOR2_X1 i_8_0_596 (.A1(n_8_0_49), .A2(n_8_0_19), .ZN(n_8_858));
   NOR2_X1 i_8_0_597 (.A1(n_8_0_49), .A2(n_8_0_20), .ZN(n_8_859));
   NOR2_X1 i_8_0_598 (.A1(n_8_0_49), .A2(n_8_0_21), .ZN(n_8_860));
   NOR2_X1 i_8_0_599 (.A1(n_8_0_49), .A2(n_8_0_22), .ZN(n_8_861));
   NOR2_X1 i_8_0_600 (.A1(n_8_0_49), .A2(n_8_0_23), .ZN(n_8_862));
   NOR2_X1 i_8_0_601 (.A1(n_8_0_49), .A2(n_8_0_24), .ZN(n_8_863));
   NOR2_X1 i_8_0_602 (.A1(n_8_0_49), .A2(n_8_0_25), .ZN(n_8_864));
   NOR2_X1 i_8_0_603 (.A1(n_8_0_49), .A2(n_8_0_26), .ZN(n_8_865));
   NOR2_X1 i_8_0_604 (.A1(n_8_0_49), .A2(n_8_0_27), .ZN(n_8_866));
   NOR2_X1 i_8_0_605 (.A1(n_8_0_49), .A2(n_8_0_28), .ZN(n_8_867));
   NOR2_X1 i_8_0_606 (.A1(n_8_0_49), .A2(n_8_0_29), .ZN(n_8_868));
   NOR2_X1 i_8_0_607 (.A1(n_8_0_49), .A2(n_8_0_30), .ZN(n_8_869));
   NOR2_X1 i_8_0_608 (.A1(n_8_0_49), .A2(n_8_0_31), .ZN(n_8_870));
   NOR2_X1 i_8_0_609 (.A1(n_8_0_49), .A2(n_8_0_32), .ZN(n_8_871));
   NOR2_X1 i_8_0_610 (.A1(n_8_0_49), .A2(n_8_0_33), .ZN(n_8_886));
   INV_X1 i_8_0_611 (.A(n_94), .ZN(n_8_0_50));
   NOR2_X1 i_8_0_612 (.A1(n_8_0_50), .A2(n_8_0_1), .ZN(n_8_791));
   NOR2_X1 i_8_0_613 (.A1(n_8_0_50), .A2(n_8_0_2), .ZN(n_8_792));
   NOR2_X1 i_8_0_614 (.A1(n_8_0_50), .A2(n_8_0_3), .ZN(n_8_793));
   NOR2_X1 i_8_0_615 (.A1(n_8_0_50), .A2(n_8_0_4), .ZN(n_8_794));
   NOR2_X1 i_8_0_616 (.A1(n_8_0_50), .A2(n_8_0_5), .ZN(n_8_795));
   NOR2_X1 i_8_0_617 (.A1(n_8_0_50), .A2(n_8_0_6), .ZN(n_8_796));
   NOR2_X1 i_8_0_618 (.A1(n_8_0_50), .A2(n_8_0_7), .ZN(n_8_797));
   NOR2_X1 i_8_0_619 (.A1(n_8_0_50), .A2(n_8_0_8), .ZN(n_8_798));
   NOR2_X1 i_8_0_620 (.A1(n_8_0_50), .A2(n_8_0_9), .ZN(n_8_799));
   NOR2_X1 i_8_0_621 (.A1(n_8_0_50), .A2(n_8_0_10), .ZN(n_8_800));
   NOR2_X1 i_8_0_622 (.A1(n_8_0_50), .A2(n_8_0_11), .ZN(n_8_801));
   NOR2_X1 i_8_0_623 (.A1(n_8_0_50), .A2(n_8_0_12), .ZN(n_8_802));
   NOR2_X1 i_8_0_624 (.A1(n_8_0_50), .A2(n_8_0_13), .ZN(n_8_803));
   NOR2_X1 i_8_0_625 (.A1(n_8_0_50), .A2(n_8_0_14), .ZN(n_8_804));
   NOR2_X1 i_8_0_626 (.A1(n_8_0_50), .A2(n_8_0_15), .ZN(n_8_805));
   NOR2_X1 i_8_0_627 (.A1(n_8_0_50), .A2(n_8_0_16), .ZN(n_8_806));
   NOR2_X1 i_8_0_628 (.A1(n_8_0_50), .A2(n_8_0_17), .ZN(n_8_807));
   NOR2_X1 i_8_0_629 (.A1(n_8_0_50), .A2(n_8_0_18), .ZN(n_8_808));
   NOR2_X1 i_8_0_630 (.A1(n_8_0_50), .A2(n_8_0_19), .ZN(n_8_809));
   NOR2_X1 i_8_0_631 (.A1(n_8_0_50), .A2(n_8_0_20), .ZN(n_8_810));
   NOR2_X1 i_8_0_632 (.A1(n_8_0_50), .A2(n_8_0_21), .ZN(n_8_811));
   NOR2_X1 i_8_0_633 (.A1(n_8_0_50), .A2(n_8_0_22), .ZN(n_8_812));
   NOR2_X1 i_8_0_634 (.A1(n_8_0_50), .A2(n_8_0_23), .ZN(n_8_813));
   NOR2_X1 i_8_0_635 (.A1(n_8_0_50), .A2(n_8_0_24), .ZN(n_8_814));
   NOR2_X1 i_8_0_636 (.A1(n_8_0_50), .A2(n_8_0_25), .ZN(n_8_815));
   NOR2_X1 i_8_0_637 (.A1(n_8_0_50), .A2(n_8_0_26), .ZN(n_8_816));
   NOR2_X1 i_8_0_638 (.A1(n_8_0_50), .A2(n_8_0_27), .ZN(n_8_817));
   NOR2_X1 i_8_0_639 (.A1(n_8_0_50), .A2(n_8_0_28), .ZN(n_8_818));
   NOR2_X1 i_8_0_640 (.A1(n_8_0_50), .A2(n_8_0_29), .ZN(n_8_819));
   NOR2_X1 i_8_0_641 (.A1(n_8_0_50), .A2(n_8_0_30), .ZN(n_8_820));
   NOR2_X1 i_8_0_642 (.A1(n_8_0_50), .A2(n_8_0_31), .ZN(n_8_821));
   NOR2_X1 i_8_0_643 (.A1(n_8_0_50), .A2(n_8_0_32), .ZN(n_8_822));
   NOR2_X1 i_8_0_644 (.A1(n_8_0_50), .A2(n_8_0_33), .ZN(n_8_838));
   INV_X1 i_8_0_645 (.A(n_125), .ZN(n_8_0_51));
   NOR2_X1 i_8_0_646 (.A1(n_8_0_51), .A2(n_8_0_1), .ZN(n_8_741));
   NOR2_X1 i_8_0_647 (.A1(n_8_0_51), .A2(n_8_0_2), .ZN(n_8_742));
   NOR2_X1 i_8_0_648 (.A1(n_8_0_51), .A2(n_8_0_3), .ZN(n_8_743));
   NOR2_X1 i_8_0_649 (.A1(n_8_0_51), .A2(n_8_0_4), .ZN(n_8_744));
   NOR2_X1 i_8_0_650 (.A1(n_8_0_51), .A2(n_8_0_5), .ZN(n_8_745));
   NOR2_X1 i_8_0_651 (.A1(n_8_0_51), .A2(n_8_0_6), .ZN(n_8_746));
   NOR2_X1 i_8_0_652 (.A1(n_8_0_51), .A2(n_8_0_7), .ZN(n_8_747));
   NOR2_X1 i_8_0_653 (.A1(n_8_0_51), .A2(n_8_0_8), .ZN(n_8_748));
   NOR2_X1 i_8_0_654 (.A1(n_8_0_51), .A2(n_8_0_9), .ZN(n_8_749));
   NOR2_X1 i_8_0_655 (.A1(n_8_0_51), .A2(n_8_0_10), .ZN(n_8_750));
   NOR2_X1 i_8_0_656 (.A1(n_8_0_51), .A2(n_8_0_11), .ZN(n_8_751));
   NOR2_X1 i_8_0_657 (.A1(n_8_0_51), .A2(n_8_0_12), .ZN(n_8_752));
   NOR2_X1 i_8_0_658 (.A1(n_8_0_51), .A2(n_8_0_13), .ZN(n_8_753));
   NOR2_X1 i_8_0_659 (.A1(n_8_0_51), .A2(n_8_0_14), .ZN(n_8_754));
   NOR2_X1 i_8_0_660 (.A1(n_8_0_51), .A2(n_8_0_15), .ZN(n_8_755));
   NOR2_X1 i_8_0_661 (.A1(n_8_0_51), .A2(n_8_0_16), .ZN(n_8_756));
   NOR2_X1 i_8_0_662 (.A1(n_8_0_51), .A2(n_8_0_17), .ZN(n_8_757));
   NOR2_X1 i_8_0_663 (.A1(n_8_0_51), .A2(n_8_0_18), .ZN(n_8_758));
   NOR2_X1 i_8_0_664 (.A1(n_8_0_51), .A2(n_8_0_19), .ZN(n_8_759));
   NOR2_X1 i_8_0_665 (.A1(n_8_0_51), .A2(n_8_0_20), .ZN(n_8_760));
   NOR2_X1 i_8_0_666 (.A1(n_8_0_51), .A2(n_8_0_21), .ZN(n_8_761));
   NOR2_X1 i_8_0_667 (.A1(n_8_0_51), .A2(n_8_0_22), .ZN(n_8_762));
   NOR2_X1 i_8_0_668 (.A1(n_8_0_51), .A2(n_8_0_23), .ZN(n_8_763));
   NOR2_X1 i_8_0_669 (.A1(n_8_0_51), .A2(n_8_0_24), .ZN(n_8_764));
   NOR2_X1 i_8_0_670 (.A1(n_8_0_51), .A2(n_8_0_25), .ZN(n_8_765));
   NOR2_X1 i_8_0_671 (.A1(n_8_0_51), .A2(n_8_0_26), .ZN(n_8_766));
   NOR2_X1 i_8_0_672 (.A1(n_8_0_51), .A2(n_8_0_27), .ZN(n_8_767));
   NOR2_X1 i_8_0_673 (.A1(n_8_0_51), .A2(n_8_0_28), .ZN(n_8_768));
   NOR2_X1 i_8_0_674 (.A1(n_8_0_51), .A2(n_8_0_29), .ZN(n_8_769));
   NOR2_X1 i_8_0_675 (.A1(n_8_0_51), .A2(n_8_0_30), .ZN(n_8_770));
   NOR2_X1 i_8_0_676 (.A1(n_8_0_51), .A2(n_8_0_31), .ZN(n_8_771));
   NOR2_X1 i_8_0_677 (.A1(n_8_0_51), .A2(n_8_0_32), .ZN(n_8_772));
   NOR2_X1 i_8_0_678 (.A1(n_8_0_51), .A2(n_8_0_33), .ZN(n_8_789));
   INV_X1 i_8_0_679 (.A(n_93), .ZN(n_8_0_52));
   NOR2_X1 i_8_0_680 (.A1(n_8_0_52), .A2(n_8_0_1), .ZN(n_8_690));
   NOR2_X1 i_8_0_681 (.A1(n_8_0_52), .A2(n_8_0_2), .ZN(n_8_691));
   NOR2_X1 i_8_0_682 (.A1(n_8_0_52), .A2(n_8_0_3), .ZN(n_8_692));
   NOR2_X1 i_8_0_683 (.A1(n_8_0_52), .A2(n_8_0_4), .ZN(n_8_693));
   NOR2_X1 i_8_0_684 (.A1(n_8_0_52), .A2(n_8_0_5), .ZN(n_8_694));
   NOR2_X1 i_8_0_685 (.A1(n_8_0_52), .A2(n_8_0_6), .ZN(n_8_695));
   NOR2_X1 i_8_0_686 (.A1(n_8_0_52), .A2(n_8_0_7), .ZN(n_8_696));
   NOR2_X1 i_8_0_687 (.A1(n_8_0_52), .A2(n_8_0_8), .ZN(n_8_697));
   NOR2_X1 i_8_0_688 (.A1(n_8_0_52), .A2(n_8_0_9), .ZN(n_8_698));
   NOR2_X1 i_8_0_689 (.A1(n_8_0_52), .A2(n_8_0_10), .ZN(n_8_699));
   NOR2_X1 i_8_0_690 (.A1(n_8_0_52), .A2(n_8_0_11), .ZN(n_8_700));
   NOR2_X1 i_8_0_691 (.A1(n_8_0_52), .A2(n_8_0_12), .ZN(n_8_701));
   NOR2_X1 i_8_0_692 (.A1(n_8_0_52), .A2(n_8_0_13), .ZN(n_8_702));
   NOR2_X1 i_8_0_693 (.A1(n_8_0_52), .A2(n_8_0_14), .ZN(n_8_703));
   NOR2_X1 i_8_0_694 (.A1(n_8_0_52), .A2(n_8_0_15), .ZN(n_8_704));
   NOR2_X1 i_8_0_695 (.A1(n_8_0_52), .A2(n_8_0_16), .ZN(n_8_705));
   NOR2_X1 i_8_0_696 (.A1(n_8_0_52), .A2(n_8_0_17), .ZN(n_8_706));
   NOR2_X1 i_8_0_697 (.A1(n_8_0_52), .A2(n_8_0_18), .ZN(n_8_707));
   NOR2_X1 i_8_0_698 (.A1(n_8_0_52), .A2(n_8_0_19), .ZN(n_8_708));
   NOR2_X1 i_8_0_699 (.A1(n_8_0_52), .A2(n_8_0_20), .ZN(n_8_709));
   NOR2_X1 i_8_0_700 (.A1(n_8_0_52), .A2(n_8_0_21), .ZN(n_8_710));
   NOR2_X1 i_8_0_701 (.A1(n_8_0_52), .A2(n_8_0_22), .ZN(n_8_711));
   NOR2_X1 i_8_0_702 (.A1(n_8_0_52), .A2(n_8_0_23), .ZN(n_8_712));
   NOR2_X1 i_8_0_703 (.A1(n_8_0_52), .A2(n_8_0_24), .ZN(n_8_713));
   NOR2_X1 i_8_0_704 (.A1(n_8_0_52), .A2(n_8_0_25), .ZN(n_8_714));
   NOR2_X1 i_8_0_705 (.A1(n_8_0_52), .A2(n_8_0_26), .ZN(n_8_715));
   NOR2_X1 i_8_0_706 (.A1(n_8_0_52), .A2(n_8_0_27), .ZN(n_8_716));
   NOR2_X1 i_8_0_707 (.A1(n_8_0_52), .A2(n_8_0_28), .ZN(n_8_717));
   NOR2_X1 i_8_0_708 (.A1(n_8_0_52), .A2(n_8_0_29), .ZN(n_8_718));
   NOR2_X1 i_8_0_709 (.A1(n_8_0_52), .A2(n_8_0_30), .ZN(n_8_719));
   NOR2_X1 i_8_0_710 (.A1(n_8_0_52), .A2(n_8_0_31), .ZN(n_8_720));
   NOR2_X1 i_8_0_711 (.A1(n_8_0_52), .A2(n_8_0_32), .ZN(n_8_721));
   NOR2_X1 i_8_0_712 (.A1(n_8_0_52), .A2(n_8_0_33), .ZN(n_8_739));
   INV_X1 i_8_0_713 (.A(n_67), .ZN(n_8_0_53));
   NOR2_X1 i_8_0_714 (.A1(n_8_0_53), .A2(n_8_0_1), .ZN(n_8_638));
   NOR2_X1 i_8_0_715 (.A1(n_8_0_53), .A2(n_8_0_2), .ZN(n_8_639));
   NOR2_X1 i_8_0_716 (.A1(n_8_0_53), .A2(n_8_0_3), .ZN(n_8_640));
   NOR2_X1 i_8_0_717 (.A1(n_8_0_53), .A2(n_8_0_4), .ZN(n_8_641));
   NOR2_X1 i_8_0_718 (.A1(n_8_0_53), .A2(n_8_0_5), .ZN(n_8_642));
   NOR2_X1 i_8_0_719 (.A1(n_8_0_53), .A2(n_8_0_6), .ZN(n_8_643));
   NOR2_X1 i_8_0_720 (.A1(n_8_0_53), .A2(n_8_0_7), .ZN(n_8_644));
   NOR2_X1 i_8_0_721 (.A1(n_8_0_53), .A2(n_8_0_8), .ZN(n_8_645));
   NOR2_X1 i_8_0_722 (.A1(n_8_0_53), .A2(n_8_0_9), .ZN(n_8_646));
   NOR2_X1 i_8_0_723 (.A1(n_8_0_53), .A2(n_8_0_10), .ZN(n_8_647));
   NOR2_X1 i_8_0_724 (.A1(n_8_0_53), .A2(n_8_0_11), .ZN(n_8_648));
   NOR2_X1 i_8_0_725 (.A1(n_8_0_53), .A2(n_8_0_12), .ZN(n_8_649));
   NOR2_X1 i_8_0_726 (.A1(n_8_0_53), .A2(n_8_0_13), .ZN(n_8_650));
   NOR2_X1 i_8_0_727 (.A1(n_8_0_53), .A2(n_8_0_14), .ZN(n_8_651));
   NOR2_X1 i_8_0_728 (.A1(n_8_0_53), .A2(n_8_0_15), .ZN(n_8_652));
   NOR2_X1 i_8_0_729 (.A1(n_8_0_53), .A2(n_8_0_16), .ZN(n_8_653));
   NOR2_X1 i_8_0_730 (.A1(n_8_0_53), .A2(n_8_0_17), .ZN(n_8_654));
   NOR2_X1 i_8_0_731 (.A1(n_8_0_53), .A2(n_8_0_18), .ZN(n_8_655));
   NOR2_X1 i_8_0_732 (.A1(n_8_0_53), .A2(n_8_0_19), .ZN(n_8_656));
   NOR2_X1 i_8_0_733 (.A1(n_8_0_53), .A2(n_8_0_20), .ZN(n_8_657));
   NOR2_X1 i_8_0_734 (.A1(n_8_0_53), .A2(n_8_0_21), .ZN(n_8_658));
   NOR2_X1 i_8_0_735 (.A1(n_8_0_53), .A2(n_8_0_22), .ZN(n_8_659));
   NOR2_X1 i_8_0_736 (.A1(n_8_0_53), .A2(n_8_0_23), .ZN(n_8_660));
   NOR2_X1 i_8_0_737 (.A1(n_8_0_53), .A2(n_8_0_24), .ZN(n_8_661));
   NOR2_X1 i_8_0_738 (.A1(n_8_0_53), .A2(n_8_0_25), .ZN(n_8_662));
   NOR2_X1 i_8_0_739 (.A1(n_8_0_53), .A2(n_8_0_26), .ZN(n_8_663));
   NOR2_X1 i_8_0_740 (.A1(n_8_0_53), .A2(n_8_0_27), .ZN(n_8_664));
   NOR2_X1 i_8_0_741 (.A1(n_8_0_53), .A2(n_8_0_28), .ZN(n_8_665));
   NOR2_X1 i_8_0_742 (.A1(n_8_0_53), .A2(n_8_0_29), .ZN(n_8_666));
   NOR2_X1 i_8_0_743 (.A1(n_8_0_53), .A2(n_8_0_30), .ZN(n_8_667));
   NOR2_X1 i_8_0_744 (.A1(n_8_0_53), .A2(n_8_0_31), .ZN(n_8_668));
   NOR2_X1 i_8_0_745 (.A1(n_8_0_53), .A2(n_8_0_32), .ZN(n_8_669));
   NOR2_X1 i_8_0_746 (.A1(n_8_0_53), .A2(n_8_0_33), .ZN(n_8_688));
   INV_X1 i_8_0_747 (.A(n_124), .ZN(n_8_0_54));
   NOR2_X1 i_8_0_748 (.A1(n_8_0_54), .A2(n_8_0_1), .ZN(n_8_585));
   NOR2_X1 i_8_0_749 (.A1(n_8_0_54), .A2(n_8_0_2), .ZN(n_8_586));
   NOR2_X1 i_8_0_750 (.A1(n_8_0_54), .A2(n_8_0_3), .ZN(n_8_587));
   NOR2_X1 i_8_0_751 (.A1(n_8_0_54), .A2(n_8_0_4), .ZN(n_8_588));
   NOR2_X1 i_8_0_752 (.A1(n_8_0_54), .A2(n_8_0_5), .ZN(n_8_589));
   NOR2_X1 i_8_0_753 (.A1(n_8_0_54), .A2(n_8_0_6), .ZN(n_8_590));
   NOR2_X1 i_8_0_754 (.A1(n_8_0_54), .A2(n_8_0_7), .ZN(n_8_591));
   NOR2_X1 i_8_0_755 (.A1(n_8_0_54), .A2(n_8_0_8), .ZN(n_8_592));
   NOR2_X1 i_8_0_756 (.A1(n_8_0_54), .A2(n_8_0_9), .ZN(n_8_593));
   NOR2_X1 i_8_0_757 (.A1(n_8_0_54), .A2(n_8_0_10), .ZN(n_8_594));
   NOR2_X1 i_8_0_758 (.A1(n_8_0_54), .A2(n_8_0_11), .ZN(n_8_595));
   NOR2_X1 i_8_0_759 (.A1(n_8_0_54), .A2(n_8_0_12), .ZN(n_8_596));
   NOR2_X1 i_8_0_760 (.A1(n_8_0_54), .A2(n_8_0_13), .ZN(n_8_597));
   NOR2_X1 i_8_0_761 (.A1(n_8_0_54), .A2(n_8_0_14), .ZN(n_8_598));
   NOR2_X1 i_8_0_762 (.A1(n_8_0_54), .A2(n_8_0_15), .ZN(n_8_599));
   NOR2_X1 i_8_0_763 (.A1(n_8_0_54), .A2(n_8_0_16), .ZN(n_8_600));
   NOR2_X1 i_8_0_764 (.A1(n_8_0_54), .A2(n_8_0_17), .ZN(n_8_601));
   NOR2_X1 i_8_0_765 (.A1(n_8_0_54), .A2(n_8_0_18), .ZN(n_8_602));
   NOR2_X1 i_8_0_766 (.A1(n_8_0_54), .A2(n_8_0_19), .ZN(n_8_603));
   NOR2_X1 i_8_0_767 (.A1(n_8_0_54), .A2(n_8_0_20), .ZN(n_8_604));
   NOR2_X1 i_8_0_768 (.A1(n_8_0_54), .A2(n_8_0_21), .ZN(n_8_605));
   NOR2_X1 i_8_0_769 (.A1(n_8_0_54), .A2(n_8_0_22), .ZN(n_8_606));
   NOR2_X1 i_8_0_770 (.A1(n_8_0_54), .A2(n_8_0_23), .ZN(n_8_607));
   NOR2_X1 i_8_0_771 (.A1(n_8_0_54), .A2(n_8_0_24), .ZN(n_8_608));
   NOR2_X1 i_8_0_772 (.A1(n_8_0_54), .A2(n_8_0_25), .ZN(n_8_609));
   NOR2_X1 i_8_0_773 (.A1(n_8_0_54), .A2(n_8_0_26), .ZN(n_8_610));
   NOR2_X1 i_8_0_774 (.A1(n_8_0_54), .A2(n_8_0_27), .ZN(n_8_611));
   NOR2_X1 i_8_0_775 (.A1(n_8_0_54), .A2(n_8_0_28), .ZN(n_8_612));
   NOR2_X1 i_8_0_776 (.A1(n_8_0_54), .A2(n_8_0_29), .ZN(n_8_613));
   NOR2_X1 i_8_0_777 (.A1(n_8_0_54), .A2(n_8_0_30), .ZN(n_8_614));
   NOR2_X1 i_8_0_778 (.A1(n_8_0_54), .A2(n_8_0_31), .ZN(n_8_615));
   NOR2_X1 i_8_0_779 (.A1(n_8_0_54), .A2(n_8_0_32), .ZN(n_8_616));
   NOR2_X1 i_8_0_780 (.A1(n_8_0_54), .A2(n_8_0_33), .ZN(n_8_636));
   INV_X1 i_8_0_781 (.A(n_92), .ZN(n_8_0_55));
   NOR2_X1 i_8_0_782 (.A1(n_8_0_55), .A2(n_8_0_1), .ZN(n_8_531));
   NOR2_X1 i_8_0_783 (.A1(n_8_0_55), .A2(n_8_0_2), .ZN(n_8_532));
   NOR2_X1 i_8_0_784 (.A1(n_8_0_55), .A2(n_8_0_3), .ZN(n_8_533));
   NOR2_X1 i_8_0_785 (.A1(n_8_0_55), .A2(n_8_0_4), .ZN(n_8_534));
   NOR2_X1 i_8_0_786 (.A1(n_8_0_55), .A2(n_8_0_5), .ZN(n_8_535));
   NOR2_X1 i_8_0_787 (.A1(n_8_0_55), .A2(n_8_0_6), .ZN(n_8_536));
   NOR2_X1 i_8_0_788 (.A1(n_8_0_55), .A2(n_8_0_7), .ZN(n_8_537));
   NOR2_X1 i_8_0_789 (.A1(n_8_0_55), .A2(n_8_0_8), .ZN(n_8_538));
   NOR2_X1 i_8_0_790 (.A1(n_8_0_55), .A2(n_8_0_9), .ZN(n_8_539));
   NOR2_X1 i_8_0_791 (.A1(n_8_0_55), .A2(n_8_0_10), .ZN(n_8_540));
   NOR2_X1 i_8_0_792 (.A1(n_8_0_55), .A2(n_8_0_11), .ZN(n_8_541));
   NOR2_X1 i_8_0_793 (.A1(n_8_0_55), .A2(n_8_0_12), .ZN(n_8_542));
   NOR2_X1 i_8_0_794 (.A1(n_8_0_55), .A2(n_8_0_13), .ZN(n_8_543));
   NOR2_X1 i_8_0_795 (.A1(n_8_0_55), .A2(n_8_0_14), .ZN(n_8_544));
   NOR2_X1 i_8_0_796 (.A1(n_8_0_55), .A2(n_8_0_15), .ZN(n_8_545));
   NOR2_X1 i_8_0_797 (.A1(n_8_0_55), .A2(n_8_0_16), .ZN(n_8_546));
   NOR2_X1 i_8_0_798 (.A1(n_8_0_55), .A2(n_8_0_17), .ZN(n_8_547));
   NOR2_X1 i_8_0_799 (.A1(n_8_0_55), .A2(n_8_0_18), .ZN(n_8_548));
   NOR2_X1 i_8_0_800 (.A1(n_8_0_55), .A2(n_8_0_19), .ZN(n_8_549));
   NOR2_X1 i_8_0_801 (.A1(n_8_0_55), .A2(n_8_0_20), .ZN(n_8_550));
   NOR2_X1 i_8_0_802 (.A1(n_8_0_55), .A2(n_8_0_21), .ZN(n_8_551));
   NOR2_X1 i_8_0_803 (.A1(n_8_0_55), .A2(n_8_0_22), .ZN(n_8_552));
   NOR2_X1 i_8_0_804 (.A1(n_8_0_55), .A2(n_8_0_23), .ZN(n_8_553));
   NOR2_X1 i_8_0_805 (.A1(n_8_0_55), .A2(n_8_0_24), .ZN(n_8_554));
   NOR2_X1 i_8_0_806 (.A1(n_8_0_55), .A2(n_8_0_25), .ZN(n_8_555));
   NOR2_X1 i_8_0_807 (.A1(n_8_0_55), .A2(n_8_0_26), .ZN(n_8_556));
   NOR2_X1 i_8_0_808 (.A1(n_8_0_55), .A2(n_8_0_27), .ZN(n_8_557));
   NOR2_X1 i_8_0_809 (.A1(n_8_0_55), .A2(n_8_0_28), .ZN(n_8_558));
   NOR2_X1 i_8_0_810 (.A1(n_8_0_55), .A2(n_8_0_29), .ZN(n_8_559));
   NOR2_X1 i_8_0_811 (.A1(n_8_0_55), .A2(n_8_0_30), .ZN(n_8_560));
   NOR2_X1 i_8_0_812 (.A1(n_8_0_55), .A2(n_8_0_31), .ZN(n_8_561));
   NOR2_X1 i_8_0_813 (.A1(n_8_0_55), .A2(n_8_0_32), .ZN(n_8_562));
   NOR2_X1 i_8_0_814 (.A1(n_8_0_55), .A2(n_8_0_33), .ZN(n_8_583));
   NOR2_X1 i_8_0_816 (.A1(n_8_0_56), .A2(n_8_0_1), .ZN(n_8_476));
   NOR2_X1 i_8_0_817 (.A1(n_8_0_56), .A2(n_8_0_2), .ZN(n_8_477));
   NOR2_X1 i_8_0_818 (.A1(n_8_0_56), .A2(n_8_0_3), .ZN(n_8_478));
   NOR2_X1 i_8_0_819 (.A1(n_8_0_56), .A2(n_8_0_4), .ZN(n_8_479));
   NOR2_X1 i_8_0_820 (.A1(n_8_0_56), .A2(n_8_0_5), .ZN(n_8_480));
   NOR2_X1 i_8_0_821 (.A1(n_8_0_56), .A2(n_8_0_6), .ZN(n_8_481));
   NOR2_X1 i_8_0_822 (.A1(n_8_0_56), .A2(n_8_0_7), .ZN(n_8_482));
   NOR2_X1 i_8_0_823 (.A1(n_8_0_56), .A2(n_8_0_8), .ZN(n_8_483));
   NOR2_X1 i_8_0_824 (.A1(n_8_0_56), .A2(n_8_0_9), .ZN(n_8_484));
   NOR2_X1 i_8_0_825 (.A1(n_8_0_56), .A2(n_8_0_10), .ZN(n_8_485));
   NOR2_X1 i_8_0_826 (.A1(n_8_0_56), .A2(n_8_0_11), .ZN(n_8_486));
   NOR2_X1 i_8_0_827 (.A1(n_8_0_56), .A2(n_8_0_12), .ZN(n_8_487));
   NOR2_X1 i_8_0_828 (.A1(n_8_0_56), .A2(n_8_0_13), .ZN(n_8_488));
   NOR2_X1 i_8_0_829 (.A1(n_8_0_56), .A2(n_8_0_14), .ZN(n_8_489));
   NOR2_X1 i_8_0_830 (.A1(n_8_0_56), .A2(n_8_0_15), .ZN(n_8_490));
   NOR2_X1 i_8_0_831 (.A1(n_8_0_56), .A2(n_8_0_16), .ZN(n_8_491));
   NOR2_X1 i_8_0_832 (.A1(n_8_0_56), .A2(n_8_0_17), .ZN(n_8_492));
   NOR2_X1 i_8_0_833 (.A1(n_8_0_56), .A2(n_8_0_18), .ZN(n_8_493));
   NOR2_X1 i_8_0_834 (.A1(n_8_0_56), .A2(n_8_0_19), .ZN(n_8_494));
   NOR2_X1 i_8_0_835 (.A1(n_8_0_56), .A2(n_8_0_20), .ZN(n_8_495));
   NOR2_X1 i_8_0_836 (.A1(n_8_0_56), .A2(n_8_0_21), .ZN(n_8_496));
   NOR2_X1 i_8_0_837 (.A1(n_8_0_56), .A2(n_8_0_22), .ZN(n_8_497));
   NOR2_X1 i_8_0_838 (.A1(n_8_0_56), .A2(n_8_0_23), .ZN(n_8_498));
   NOR2_X1 i_8_0_839 (.A1(n_8_0_56), .A2(n_8_0_24), .ZN(n_8_499));
   NOR2_X1 i_8_0_840 (.A1(n_8_0_56), .A2(n_8_0_25), .ZN(n_8_500));
   NOR2_X1 i_8_0_841 (.A1(n_8_0_56), .A2(n_8_0_26), .ZN(n_8_501));
   NOR2_X1 i_8_0_842 (.A1(n_8_0_56), .A2(n_8_0_27), .ZN(n_8_502));
   NOR2_X1 i_8_0_843 (.A1(n_8_0_56), .A2(n_8_0_28), .ZN(n_8_503));
   NOR2_X1 i_8_0_844 (.A1(n_8_0_56), .A2(n_8_0_29), .ZN(n_8_504));
   NOR2_X1 i_8_0_846 (.A1(n_8_0_56), .A2(n_8_0_31), .ZN(n_8_506));
   NOR2_X1 i_8_0_847 (.A1(n_8_0_56), .A2(n_8_0_32), .ZN(n_8_507));
   NOR2_X1 i_8_0_848 (.A1(n_8_0_56), .A2(n_8_0_33), .ZN(n_8_526));
   NOR2_X1 i_8_0_850 (.A1(n_8_0_57), .A2(n_8_0_1), .ZN(n_8_420));
   NOR2_X1 i_8_0_851 (.A1(n_8_0_57), .A2(n_8_0_2), .ZN(n_8_421));
   NOR2_X1 i_8_0_852 (.A1(n_8_0_57), .A2(n_8_0_3), .ZN(n_8_422));
   NOR2_X1 i_8_0_853 (.A1(n_8_0_57), .A2(n_8_0_4), .ZN(n_8_423));
   NOR2_X1 i_8_0_854 (.A1(n_8_0_57), .A2(n_8_0_5), .ZN(n_8_424));
   NOR2_X1 i_8_0_855 (.A1(n_8_0_57), .A2(n_8_0_6), .ZN(n_8_425));
   NOR2_X1 i_8_0_856 (.A1(n_8_0_57), .A2(n_8_0_7), .ZN(n_8_426));
   NOR2_X1 i_8_0_857 (.A1(n_8_0_57), .A2(n_8_0_8), .ZN(n_8_427));
   NOR2_X1 i_8_0_858 (.A1(n_8_0_57), .A2(n_8_0_9), .ZN(n_8_428));
   NOR2_X1 i_8_0_859 (.A1(n_8_0_57), .A2(n_8_0_10), .ZN(n_8_429));
   NOR2_X1 i_8_0_860 (.A1(n_8_0_57), .A2(n_8_0_11), .ZN(n_8_430));
   NOR2_X1 i_8_0_861 (.A1(n_8_0_57), .A2(n_8_0_12), .ZN(n_8_431));
   NOR2_X1 i_8_0_862 (.A1(n_8_0_57), .A2(n_8_0_13), .ZN(n_8_432));
   NOR2_X1 i_8_0_863 (.A1(n_8_0_57), .A2(n_8_0_14), .ZN(n_8_433));
   NOR2_X1 i_8_0_864 (.A1(n_8_0_57), .A2(n_8_0_15), .ZN(n_8_434));
   NOR2_X1 i_8_0_865 (.A1(n_8_0_57), .A2(n_8_0_16), .ZN(n_8_435));
   NOR2_X1 i_8_0_866 (.A1(n_8_0_57), .A2(n_8_0_17), .ZN(n_8_436));
   NOR2_X1 i_8_0_867 (.A1(n_8_0_57), .A2(n_8_0_18), .ZN(n_8_437));
   NOR2_X1 i_8_0_868 (.A1(n_8_0_57), .A2(n_8_0_19), .ZN(n_8_438));
   NOR2_X1 i_8_0_869 (.A1(n_8_0_57), .A2(n_8_0_20), .ZN(n_8_439));
   NOR2_X1 i_8_0_870 (.A1(n_8_0_57), .A2(n_8_0_21), .ZN(n_8_440));
   NOR2_X1 i_8_0_871 (.A1(n_8_0_57), .A2(n_8_0_22), .ZN(n_8_441));
   NOR2_X1 i_8_0_872 (.A1(n_8_0_57), .A2(n_8_0_23), .ZN(n_8_442));
   NOR2_X1 i_8_0_873 (.A1(n_8_0_57), .A2(n_8_0_24), .ZN(n_8_443));
   NOR2_X1 i_8_0_874 (.A1(n_8_0_57), .A2(n_8_0_25), .ZN(n_8_444));
   NOR2_X1 i_8_0_875 (.A1(n_8_0_57), .A2(n_8_0_26), .ZN(n_8_445));
   NOR2_X1 i_8_0_876 (.A1(n_8_0_57), .A2(n_8_0_27), .ZN(n_8_446));
   NOR2_X1 i_8_0_877 (.A1(n_8_0_57), .A2(n_8_0_28), .ZN(n_8_447));
   NOR2_X1 i_8_0_879 (.A1(n_8_0_57), .A2(n_8_0_30), .ZN(n_8_449));
   NOR2_X1 i_8_0_881 (.A1(n_8_0_57), .A2(n_8_0_32), .ZN(n_8_451));
   NOR2_X1 i_8_0_882 (.A1(n_8_0_57), .A2(n_8_0_33), .ZN(n_8_471));
   NOR2_X1 i_8_0_884 (.A1(n_8_0_58), .A2(n_8_0_1), .ZN(n_8_399));
   NOR2_X1 i_8_0_885 (.A1(n_8_0_58), .A2(n_8_0_2), .ZN(n_8_400));
   NOR2_X1 i_8_0_886 (.A1(n_8_0_58), .A2(n_8_0_3), .ZN(n_8_401));
   NOR2_X1 i_8_0_887 (.A1(n_8_0_58), .A2(n_8_0_4), .ZN(n_8_402));
   NOR2_X1 i_8_0_888 (.A1(n_8_0_58), .A2(n_8_0_5), .ZN(n_8_403));
   NOR2_X1 i_8_0_889 (.A1(n_8_0_58), .A2(n_8_0_6), .ZN(n_8_404));
   NOR2_X1 i_8_0_890 (.A1(n_8_0_58), .A2(n_8_0_7), .ZN(n_8_405));
   NOR2_X1 i_8_0_891 (.A1(n_8_0_58), .A2(n_8_0_8), .ZN(n_8_406));
   NOR2_X1 i_8_0_892 (.A1(n_8_0_58), .A2(n_8_0_9), .ZN(n_8_407));
   NOR2_X1 i_8_0_893 (.A1(n_8_0_58), .A2(n_8_0_10), .ZN(n_8_408));
   NOR2_X1 i_8_0_894 (.A1(n_8_0_58), .A2(n_8_0_11), .ZN(n_8_409));
   NOR2_X1 i_8_0_895 (.A1(n_8_0_58), .A2(n_8_0_12), .ZN(n_8_410));
   NOR2_X1 i_8_0_896 (.A1(n_8_0_58), .A2(n_8_0_13), .ZN(n_8_411));
   NOR2_X1 i_8_0_897 (.A1(n_8_0_58), .A2(n_8_0_14), .ZN(n_8_412));
   NOR2_X1 i_8_0_898 (.A1(n_8_0_58), .A2(n_8_0_15), .ZN(n_8_413));
   NOR2_X1 i_8_0_899 (.A1(n_8_0_58), .A2(n_8_0_16), .ZN(n_8_414));
   NOR2_X1 i_8_0_900 (.A1(n_8_0_58), .A2(n_8_0_17), .ZN(n_8_415));
   NOR2_X1 i_8_0_901 (.A1(n_8_0_58), .A2(n_8_0_18), .ZN(n_8_416));
   NOR2_X1 i_8_0_902 (.A1(n_8_0_58), .A2(n_8_0_19), .ZN(n_8_417));
   NOR2_X1 i_8_0_903 (.A1(n_8_0_58), .A2(n_8_0_20), .ZN(n_8_418));
   NOR2_X1 i_8_0_904 (.A1(n_8_0_58), .A2(n_8_0_21), .ZN(n_8_419));
   NOR2_X1 i_8_0_905 (.A1(n_8_0_58), .A2(n_8_0_22), .ZN(n_8_452));
   NOR2_X1 i_8_0_906 (.A1(n_8_0_58), .A2(n_8_0_23), .ZN(n_8_453));
   NOR2_X1 i_8_0_907 (.A1(n_8_0_58), .A2(n_8_0_24), .ZN(n_8_454));
   NOR2_X1 i_8_0_908 (.A1(n_8_0_58), .A2(n_8_0_25), .ZN(n_8_455));
   NOR2_X1 i_8_0_909 (.A1(n_8_0_58), .A2(n_8_0_26), .ZN(n_8_456));
   NOR2_X1 i_8_0_910 (.A1(n_8_0_58), .A2(n_8_0_27), .ZN(n_8_457));
   NOR2_X1 i_8_0_911 (.A1(n_8_0_58), .A2(n_8_0_28), .ZN(n_8_458));
   NOR2_X1 i_8_0_912 (.A1(n_8_0_58), .A2(n_8_0_29), .ZN(n_8_459));
   NOR2_X1 i_8_0_914 (.A1(n_8_0_58), .A2(n_8_0_31), .ZN(n_8_461));
   NOR2_X1 i_8_0_916 (.A1(n_8_0_58), .A2(n_8_0_33), .ZN(n_8_463));
   NOR2_X1 i_8_0_918 (.A1(n_8_0_59), .A2(n_8_0_1), .ZN(n_8_464));
   NOR2_X1 i_8_0_919 (.A1(n_8_0_59), .A2(n_8_0_2), .ZN(n_8_465));
   NOR2_X1 i_8_0_920 (.A1(n_8_0_59), .A2(n_8_0_3), .ZN(n_8_466));
   NOR2_X1 i_8_0_921 (.A1(n_8_0_59), .A2(n_8_0_4), .ZN(n_8_467));
   NOR2_X1 i_8_0_922 (.A1(n_8_0_59), .A2(n_8_0_5), .ZN(n_8_468));
   NOR2_X1 i_8_0_923 (.A1(n_8_0_59), .A2(n_8_0_6), .ZN(n_8_469));
   NOR2_X1 i_8_0_924 (.A1(n_8_0_59), .A2(n_8_0_7), .ZN(n_8_470));
   NOR2_X1 i_8_0_925 (.A1(n_8_0_59), .A2(n_8_0_8), .ZN(n_8_472));
   NOR2_X1 i_8_0_926 (.A1(n_8_0_59), .A2(n_8_0_9), .ZN(n_8_473));
   NOR2_X1 i_8_0_927 (.A1(n_8_0_59), .A2(n_8_0_10), .ZN(n_8_474));
   NOR2_X1 i_8_0_928 (.A1(n_8_0_59), .A2(n_8_0_11), .ZN(n_8_475));
   NOR2_X1 i_8_0_929 (.A1(n_8_0_59), .A2(n_8_0_12), .ZN(n_8_508));
   NOR2_X1 i_8_0_930 (.A1(n_8_0_59), .A2(n_8_0_13), .ZN(n_8_509));
   NOR2_X1 i_8_0_931 (.A1(n_8_0_59), .A2(n_8_0_14), .ZN(n_8_510));
   NOR2_X1 i_8_0_932 (.A1(n_8_0_59), .A2(n_8_0_15), .ZN(n_8_511));
   NOR2_X1 i_8_0_933 (.A1(n_8_0_59), .A2(n_8_0_16), .ZN(n_8_512));
   NOR2_X1 i_8_0_934 (.A1(n_8_0_59), .A2(n_8_0_17), .ZN(n_8_513));
   NOR2_X1 i_8_0_935 (.A1(n_8_0_59), .A2(n_8_0_18), .ZN(n_8_514));
   NOR2_X1 i_8_0_936 (.A1(n_8_0_59), .A2(n_8_0_19), .ZN(n_8_515));
   NOR2_X1 i_8_0_937 (.A1(n_8_0_59), .A2(n_8_0_20), .ZN(n_8_516));
   NOR2_X1 i_8_0_938 (.A1(n_8_0_59), .A2(n_8_0_21), .ZN(n_8_517));
   NOR2_X1 i_8_0_939 (.A1(n_8_0_59), .A2(n_8_0_22), .ZN(n_8_518));
   NOR2_X1 i_8_0_940 (.A1(n_8_0_59), .A2(n_8_0_23), .ZN(n_8_519));
   NOR2_X1 i_8_0_941 (.A1(n_8_0_59), .A2(n_8_0_24), .ZN(n_8_520));
   NOR2_X1 i_8_0_942 (.A1(n_8_0_59), .A2(n_8_0_25), .ZN(n_8_521));
   NOR2_X1 i_8_0_943 (.A1(n_8_0_59), .A2(n_8_0_26), .ZN(n_8_522));
   NOR2_X1 i_8_0_944 (.A1(n_8_0_59), .A2(n_8_0_27), .ZN(n_8_523));
   NOR2_X1 i_8_0_945 (.A1(n_8_0_59), .A2(n_8_0_28), .ZN(n_8_524));
   NOR2_X1 i_8_0_946 (.A1(n_8_0_59), .A2(n_8_0_29), .ZN(n_8_525));
   NOR2_X1 i_8_0_949 (.A1(n_8_0_59), .A2(n_8_0_32), .ZN(n_8_529));
   NOR2_X1 i_8_0_952 (.A1(n_8_0_60), .A2(n_8_0_1), .ZN(n_8_563));
   NOR2_X1 i_8_0_953 (.A1(n_8_0_60), .A2(n_8_0_2), .ZN(n_8_564));
   NOR2_X1 i_8_0_954 (.A1(n_8_0_60), .A2(n_8_0_3), .ZN(n_8_565));
   NOR2_X1 i_8_0_955 (.A1(n_8_0_60), .A2(n_8_0_4), .ZN(n_8_566));
   NOR2_X1 i_8_0_956 (.A1(n_8_0_60), .A2(n_8_0_5), .ZN(n_8_567));
   NOR2_X1 i_8_0_957 (.A1(n_8_0_60), .A2(n_8_0_6), .ZN(n_8_568));
   NOR2_X1 i_8_0_958 (.A1(n_8_0_60), .A2(n_8_0_7), .ZN(n_8_569));
   NOR2_X1 i_8_0_959 (.A1(n_8_0_60), .A2(n_8_0_8), .ZN(n_8_570));
   NOR2_X1 i_8_0_960 (.A1(n_8_0_60), .A2(n_8_0_9), .ZN(n_8_571));
   NOR2_X1 i_8_0_961 (.A1(n_8_0_60), .A2(n_8_0_10), .ZN(n_8_572));
   NOR2_X1 i_8_0_962 (.A1(n_8_0_60), .A2(n_8_0_11), .ZN(n_8_573));
   NOR2_X1 i_8_0_963 (.A1(n_8_0_60), .A2(n_8_0_12), .ZN(n_8_574));
   NOR2_X1 i_8_0_964 (.A1(n_8_0_60), .A2(n_8_0_13), .ZN(n_8_575));
   NOR2_X1 i_8_0_965 (.A1(n_8_0_60), .A2(n_8_0_14), .ZN(n_8_576));
   NOR2_X1 i_8_0_966 (.A1(n_8_0_60), .A2(n_8_0_15), .ZN(n_8_577));
   NOR2_X1 i_8_0_967 (.A1(n_8_0_60), .A2(n_8_0_16), .ZN(n_8_578));
   NOR2_X1 i_8_0_968 (.A1(n_8_0_60), .A2(n_8_0_17), .ZN(n_8_579));
   NOR2_X1 i_8_0_969 (.A1(n_8_0_60), .A2(n_8_0_18), .ZN(n_8_580));
   NOR2_X1 i_8_0_970 (.A1(n_8_0_60), .A2(n_8_0_19), .ZN(n_8_581));
   NOR2_X1 i_8_0_971 (.A1(n_8_0_60), .A2(n_8_0_20), .ZN(n_8_582));
   NOR2_X1 i_8_0_972 (.A1(n_8_0_60), .A2(n_8_0_21), .ZN(n_8_584));
   NOR2_X1 i_8_0_973 (.A1(n_8_0_60), .A2(n_8_0_22), .ZN(n_8_617));
   NOR2_X1 i_8_0_974 (.A1(n_8_0_60), .A2(n_8_0_23), .ZN(n_8_618));
   NOR2_X1 i_8_0_975 (.A1(n_8_0_60), .A2(n_8_0_24), .ZN(n_8_619));
   NOR2_X1 i_8_0_976 (.A1(n_8_0_60), .A2(n_8_0_25), .ZN(n_8_620));
   NOR2_X1 i_8_0_977 (.A1(n_8_0_60), .A2(n_8_0_26), .ZN(n_8_621));
   NOR2_X1 i_8_0_978 (.A1(n_8_0_60), .A2(n_8_0_27), .ZN(n_8_622));
   NOR2_X1 i_8_0_979 (.A1(n_8_0_60), .A2(n_8_0_28), .ZN(n_8_623));
   NOR2_X1 i_8_0_980 (.A1(n_8_0_60), .A2(n_8_0_29), .ZN(n_8_624));
   NOR2_X1 i_8_0_981 (.A1(n_8_0_60), .A2(n_8_0_30), .ZN(n_8_625));
   NOR2_X1 i_8_0_982 (.A1(n_8_0_60), .A2(n_8_0_31), .ZN(n_8_626));
   NOR2_X1 i_8_0_986 (.A1(n_8_0_61), .A2(n_8_0_1), .ZN(n_8_629));
   NOR2_X1 i_8_0_987 (.A1(n_8_0_61), .A2(n_8_0_2), .ZN(n_8_630));
   NOR2_X1 i_8_0_988 (.A1(n_8_0_61), .A2(n_8_0_3), .ZN(n_8_631));
   NOR2_X1 i_8_0_989 (.A1(n_8_0_61), .A2(n_8_0_4), .ZN(n_8_632));
   NOR2_X1 i_8_0_990 (.A1(n_8_0_61), .A2(n_8_0_5), .ZN(n_8_633));
   NOR2_X1 i_8_0_991 (.A1(n_8_0_61), .A2(n_8_0_6), .ZN(n_8_634));
   NOR2_X1 i_8_0_992 (.A1(n_8_0_61), .A2(n_8_0_7), .ZN(n_8_635));
   NOR2_X1 i_8_0_993 (.A1(n_8_0_61), .A2(n_8_0_8), .ZN(n_8_637));
   NOR2_X1 i_8_0_994 (.A1(n_8_0_61), .A2(n_8_0_9), .ZN(n_8_670));
   NOR2_X1 i_8_0_995 (.A1(n_8_0_61), .A2(n_8_0_10), .ZN(n_8_671));
   NOR2_X1 i_8_0_996 (.A1(n_8_0_61), .A2(n_8_0_11), .ZN(n_8_672));
   NOR2_X1 i_8_0_997 (.A1(n_8_0_61), .A2(n_8_0_12), .ZN(n_8_673));
   NOR2_X1 i_8_0_998 (.A1(n_8_0_61), .A2(n_8_0_13), .ZN(n_8_674));
   NOR2_X1 i_8_0_999 (.A1(n_8_0_61), .A2(n_8_0_14), .ZN(n_8_675));
   NOR2_X1 i_8_0_1000 (.A1(n_8_0_61), .A2(n_8_0_15), .ZN(n_8_676));
   NOR2_X1 i_8_0_1001 (.A1(n_8_0_61), .A2(n_8_0_16), .ZN(n_8_677));
   NOR2_X1 i_8_0_1002 (.A1(n_8_0_61), .A2(n_8_0_17), .ZN(n_8_678));
   NOR2_X1 i_8_0_1003 (.A1(n_8_0_61), .A2(n_8_0_18), .ZN(n_8_679));
   NOR2_X1 i_8_0_1004 (.A1(n_8_0_61), .A2(n_8_0_19), .ZN(n_8_680));
   NOR2_X1 i_8_0_1005 (.A1(n_8_0_61), .A2(n_8_0_20), .ZN(n_8_681));
   NOR2_X1 i_8_0_1006 (.A1(n_8_0_61), .A2(n_8_0_21), .ZN(n_8_682));
   NOR2_X1 i_8_0_1007 (.A1(n_8_0_61), .A2(n_8_0_22), .ZN(n_8_683));
   NOR2_X1 i_8_0_1008 (.A1(n_8_0_61), .A2(n_8_0_23), .ZN(n_8_684));
   NOR2_X1 i_8_0_1009 (.A1(n_8_0_61), .A2(n_8_0_24), .ZN(n_8_685));
   NOR2_X1 i_8_0_1011 (.A1(n_8_0_61), .A2(n_8_0_26), .ZN(n_8_687));
   NOR2_X1 i_8_0_1012 (.A1(n_8_0_61), .A2(n_8_0_27), .ZN(n_8_689));
   NOR2_X1 i_8_0_1013 (.A1(n_8_0_61), .A2(n_8_0_28), .ZN(n_8_722));
   NOR2_X1 i_8_0_1014 (.A1(n_8_0_61), .A2(n_8_0_29), .ZN(n_8_723));
   NOR2_X1 i_8_0_1016 (.A1(n_8_0_61), .A2(n_8_0_31), .ZN(n_8_725));
   NOR2_X1 i_8_0_1017 (.A1(n_8_0_61), .A2(n_8_0_32), .ZN(n_8_726));
   NOR2_X1 i_8_0_1020 (.A1(n_8_0_62), .A2(n_8_0_1), .ZN(n_8_728));
   NOR2_X1 i_8_0_1021 (.A1(n_8_0_62), .A2(n_8_0_2), .ZN(n_8_729));
   NOR2_X1 i_8_0_1022 (.A1(n_8_0_62), .A2(n_8_0_3), .ZN(n_8_730));
   NOR2_X1 i_8_0_1023 (.A1(n_8_0_62), .A2(n_8_0_4), .ZN(n_8_731));
   NOR2_X1 i_8_0_1024 (.A1(n_8_0_62), .A2(n_8_0_5), .ZN(n_8_732));
   NOR2_X1 i_8_0_1025 (.A1(n_8_0_62), .A2(n_8_0_6), .ZN(n_8_733));
   NOR2_X1 i_8_0_1026 (.A1(n_8_0_62), .A2(n_8_0_7), .ZN(n_8_734));
   NOR2_X1 i_8_0_1027 (.A1(n_8_0_62), .A2(n_8_0_8), .ZN(n_8_735));
   NOR2_X1 i_8_0_1028 (.A1(n_8_0_62), .A2(n_8_0_9), .ZN(n_8_736));
   NOR2_X1 i_8_0_1029 (.A1(n_8_0_62), .A2(n_8_0_10), .ZN(n_8_737));
   NOR2_X1 i_8_0_1030 (.A1(n_8_0_62), .A2(n_8_0_11), .ZN(n_8_738));
   NOR2_X1 i_8_0_1031 (.A1(n_8_0_62), .A2(n_8_0_12), .ZN(n_8_740));
   NOR2_X1 i_8_0_1032 (.A1(n_8_0_62), .A2(n_8_0_13), .ZN(n_8_773));
   NOR2_X1 i_8_0_1033 (.A1(n_8_0_62), .A2(n_8_0_14), .ZN(n_8_774));
   NOR2_X1 i_8_0_1034 (.A1(n_8_0_62), .A2(n_8_0_15), .ZN(n_8_775));
   NOR2_X1 i_8_0_1035 (.A1(n_8_0_62), .A2(n_8_0_16), .ZN(n_8_776));
   NOR2_X1 i_8_0_1036 (.A1(n_8_0_62), .A2(n_8_0_17), .ZN(n_8_777));
   NOR2_X1 i_8_0_1037 (.A1(n_8_0_62), .A2(n_8_0_18), .ZN(n_8_778));
   NOR2_X1 i_8_0_1038 (.A1(n_8_0_62), .A2(n_8_0_19), .ZN(n_8_779));
   NOR2_X1 i_8_0_1039 (.A1(n_8_0_62), .A2(n_8_0_20), .ZN(n_8_780));
   NOR2_X1 i_8_0_1040 (.A1(n_8_0_62), .A2(n_8_0_21), .ZN(n_8_781));
   NOR2_X1 i_8_0_1041 (.A1(n_8_0_62), .A2(n_8_0_22), .ZN(n_8_782));
   NOR2_X1 i_8_0_1042 (.A1(n_8_0_62), .A2(n_8_0_23), .ZN(n_8_783));
   NOR2_X1 i_8_0_1043 (.A1(n_8_0_62), .A2(n_8_0_24), .ZN(n_8_784));
   NOR2_X1 i_8_0_1044 (.A1(n_8_0_62), .A2(n_8_0_25), .ZN(n_8_785));
   NOR2_X1 i_8_0_1046 (.A1(n_8_0_62), .A2(n_8_0_27), .ZN(n_8_787));
   NOR2_X1 i_8_0_1047 (.A1(n_8_0_62), .A2(n_8_0_28), .ZN(n_8_788));
   NOR2_X1 i_8_0_1048 (.A1(n_8_0_62), .A2(n_8_0_29), .ZN(n_8_790));
   NOR2_X1 i_8_0_1050 (.A1(n_8_0_62), .A2(n_8_0_31), .ZN(n_8_824));
   NOR2_X1 i_8_0_1051 (.A1(n_8_0_62), .A2(n_8_0_32), .ZN(n_8_825));
   NOR2_X1 i_8_0_1052 (.A1(n_8_0_62), .A2(n_8_0_33), .ZN(n_8_826));
   NOR2_X1 i_8_0_1054 (.A1(n_8_0_63), .A2(n_8_0_1), .ZN(n_8_827));
   NOR2_X1 i_8_0_1055 (.A1(n_8_0_63), .A2(n_8_0_2), .ZN(n_8_828));
   NOR2_X1 i_8_0_1056 (.A1(n_8_0_63), .A2(n_8_0_3), .ZN(n_8_829));
   NOR2_X1 i_8_0_1057 (.A1(n_8_0_63), .A2(n_8_0_4), .ZN(n_8_830));
   NOR2_X1 i_8_0_1058 (.A1(n_8_0_63), .A2(n_8_0_5), .ZN(n_8_831));
   NOR2_X1 i_8_0_1059 (.A1(n_8_0_63), .A2(n_8_0_6), .ZN(n_8_832));
   NOR2_X1 i_8_0_1060 (.A1(n_8_0_63), .A2(n_8_0_7), .ZN(n_8_833));
   NOR2_X1 i_8_0_1061 (.A1(n_8_0_63), .A2(n_8_0_8), .ZN(n_8_834));
   NOR2_X1 i_8_0_1062 (.A1(n_8_0_63), .A2(n_8_0_9), .ZN(n_8_835));
   NOR2_X1 i_8_0_1063 (.A1(n_8_0_63), .A2(n_8_0_10), .ZN(n_8_836));
   NOR2_X1 i_8_0_1064 (.A1(n_8_0_63), .A2(n_8_0_11), .ZN(n_8_837));
   NOR2_X1 i_8_0_1065 (.A1(n_8_0_63), .A2(n_8_0_12), .ZN(n_8_839));
   NOR2_X1 i_8_0_1066 (.A1(n_8_0_63), .A2(n_8_0_13), .ZN(n_8_872));
   NOR2_X1 i_8_0_1067 (.A1(n_8_0_63), .A2(n_8_0_14), .ZN(n_8_873));
   NOR2_X1 i_8_0_1068 (.A1(n_8_0_63), .A2(n_8_0_15), .ZN(n_8_874));
   NOR2_X1 i_8_0_1069 (.A1(n_8_0_63), .A2(n_8_0_16), .ZN(n_8_875));
   NOR2_X1 i_8_0_1070 (.A1(n_8_0_63), .A2(n_8_0_17), .ZN(n_8_876));
   NOR2_X1 i_8_0_1071 (.A1(n_8_0_63), .A2(n_8_0_18), .ZN(n_8_877));
   NOR2_X1 i_8_0_1072 (.A1(n_8_0_63), .A2(n_8_0_19), .ZN(n_8_878));
   NOR2_X1 i_8_0_1073 (.A1(n_8_0_63), .A2(n_8_0_20), .ZN(n_8_879));
   NOR2_X1 i_8_0_1074 (.A1(n_8_0_63), .A2(n_8_0_21), .ZN(n_8_880));
   NOR2_X1 i_8_0_1075 (.A1(n_8_0_63), .A2(n_8_0_22), .ZN(n_8_881));
   NOR2_X1 i_8_0_1076 (.A1(n_8_0_63), .A2(n_8_0_23), .ZN(n_8_882));
   NOR2_X1 i_8_0_1077 (.A1(n_8_0_63), .A2(n_8_0_24), .ZN(n_8_883));
   NOR2_X1 i_8_0_1078 (.A1(n_8_0_63), .A2(n_8_0_25), .ZN(n_8_884));
   NOR2_X1 i_8_0_1079 (.A1(n_8_0_63), .A2(n_8_0_26), .ZN(n_8_885));
   NOR2_X1 i_8_0_1081 (.A1(n_8_0_63), .A2(n_8_0_28), .ZN(n_8_920));
   NOR2_X1 i_8_0_1083 (.A1(n_8_0_63), .A2(n_8_0_30), .ZN(n_8_922));
   NOR2_X1 i_8_0_1084 (.A1(n_8_0_63), .A2(n_8_0_31), .ZN(n_8_923));
   NOR2_X1 i_8_0_1085 (.A1(n_8_0_63), .A2(n_8_0_32), .ZN(n_8_924));
   NOR2_X1 i_8_0_1086 (.A1(n_8_0_63), .A2(n_8_0_33), .ZN(n_8_925));
   NOR2_X1 i_8_0_1088 (.A1(n_8_0_1), .A2(n_8_0_64), .ZN(n_8_926));
   NOR2_X1 i_8_0_1089 (.A1(n_8_0_2), .A2(n_8_0_64), .ZN(n_8_927));
   NOR2_X1 i_8_0_1090 (.A1(n_8_0_3), .A2(n_8_0_64), .ZN(n_8_928));
   NOR2_X1 i_8_0_1091 (.A1(n_8_0_4), .A2(n_8_0_64), .ZN(n_8_929));
   NOR2_X1 i_8_0_1092 (.A1(n_8_0_5), .A2(n_8_0_64), .ZN(n_8_930));
   NOR2_X1 i_8_0_1093 (.A1(n_8_0_6), .A2(n_8_0_64), .ZN(n_8_931));
   NOR2_X1 i_8_0_1094 (.A1(n_8_0_7), .A2(n_8_0_64), .ZN(n_8_932));
   NOR2_X1 i_8_0_1095 (.A1(n_8_0_8), .A2(n_8_0_64), .ZN(n_8_934));
   NOR2_X1 i_8_0_1096 (.A1(n_8_0_9), .A2(n_8_0_64), .ZN(n_8_967));
   NOR2_X1 i_8_0_1097 (.A1(n_8_0_10), .A2(n_8_0_64), .ZN(n_8_968));
   NOR2_X1 i_8_0_1098 (.A1(n_8_0_11), .A2(n_8_0_64), .ZN(n_8_969));
   NOR2_X1 i_8_0_1099 (.A1(n_8_0_12), .A2(n_8_0_64), .ZN(n_8_970));
   NOR2_X1 i_8_0_1100 (.A1(n_8_0_13), .A2(n_8_0_64), .ZN(n_8_971));
   NOR2_X1 i_8_0_1101 (.A1(n_8_0_14), .A2(n_8_0_64), .ZN(n_8_972));
   NOR2_X1 i_8_0_1102 (.A1(n_8_0_15), .A2(n_8_0_64), .ZN(n_8_973));
   NOR2_X1 i_8_0_1103 (.A1(n_8_0_16), .A2(n_8_0_64), .ZN(n_8_974));
   NOR2_X1 i_8_0_1104 (.A1(n_8_0_17), .A2(n_8_0_64), .ZN(n_8_975));
   NOR2_X1 i_8_0_1105 (.A1(n_8_0_18), .A2(n_8_0_64), .ZN(n_8_976));
   NOR2_X1 i_8_0_1106 (.A1(n_8_0_19), .A2(n_8_0_64), .ZN(n_8_977));
   NOR2_X1 i_8_0_1107 (.A1(n_8_0_20), .A2(n_8_0_64), .ZN(n_8_978));
   NOR2_X1 i_8_0_1108 (.A1(n_8_0_21), .A2(n_8_0_64), .ZN(n_8_980));
   NOR2_X1 i_8_0_1109 (.A1(n_8_0_22), .A2(n_8_0_64), .ZN(n_8_1013));
   NOR2_X1 i_8_0_1110 (.A1(n_8_0_23), .A2(n_8_0_64), .ZN(n_8_1014));
   NOR2_X1 i_8_0_1111 (.A1(n_8_0_24), .A2(n_8_0_64), .ZN(n_8_1015));
   NOR2_X1 i_8_0_1112 (.A1(n_8_0_25), .A2(n_8_0_64), .ZN(n_8_1016));
   NOR2_X1 i_8_0_1113 (.A1(n_8_0_26), .A2(n_8_0_64), .ZN(n_8_1017));
   NOR2_X1 i_8_0_1114 (.A1(n_8_0_27), .A2(n_8_0_64), .ZN(n_8_1018));
   NOR2_X1 i_8_0_1116 (.A1(n_8_0_29), .A2(n_8_0_64), .ZN(n_8_1020));
   NOR2_X1 i_8_0_1118 (.A1(n_8_0_31), .A2(n_8_0_64), .ZN(n_8_1022));
   NOR2_X1 i_8_0_1119 (.A1(n_8_0_32), .A2(n_8_0_64), .ZN(n_8_1023));
   NOR2_X1 i_8_0_1120 (.A1(n_8_0_33), .A2(n_8_0_64), .ZN(n_8_1025));
   INV_X1 i_8_0_0 (.A(n_64), .ZN(n_8_0_65));
   INV_X1 i_8_0_1 (.A(n_65), .ZN(n_8_0_66));
   INV_X1 i_8_0_3 (.A(n_66), .ZN(n_8_0_67));
   INV_X1 i_8_0_5 (.A(n_87), .ZN(n_8_0_68));
   INV_X1 i_8_0_7 (.A(n_88), .ZN(n_8_0_69));
   INV_X1 i_8_0_9 (.A(n_89), .ZN(n_8_0_70));
   INV_X1 i_8_0_13 (.A(n_90), .ZN(n_8_0_71));
   INV_X1 i_8_0_17 (.A(n_91), .ZN(n_8_0_72));
   INV_X1 i_8_0_21 (.A(n_103), .ZN(n_8_0_73));
   INV_X1 i_8_0_23 (.A(n_104), .ZN(n_8_0_74));
   INV_X1 i_8_0_25 (.A(n_105), .ZN(n_8_0_75));
   INV_X1 i_8_0_49 (.A(n_79), .ZN(n_8_0_76));
   INV_X1 i_8_0_51 (.A(n_80), .ZN(n_8_0_77));
   INV_X1 i_8_0_53 (.A(n_81), .ZN(n_8_0_78));
   INV_X1 i_8_0_54 (.A(n_77), .ZN(n_8_0_79));
   INV_X1 i_8_0_55 (.A(n_75), .ZN(n_8_0_80));
   INV_X1 i_8_0_57 (.A(n_85), .ZN(n_8_0_81));
   INV_X1 i_8_0_58 (.A(n_74), .ZN(n_8_0_82));
   INV_X1 i_8_0_59 (.A(n_123), .ZN(n_8_0_83));
   INV_X1 i_8_0_60 (.A(n_122), .ZN(n_8_0_84));
   INV_X1 i_8_0_61 (.A(n_73), .ZN(n_8_0_85));
   INV_X1 i_8_0_63 (.A(n_84), .ZN(n_8_0_86));
   INV_X1 i_8_0_65 (.A(n_114), .ZN(n_8_0_87));
   INV_X1 i_8_0_101 (.A(n_113), .ZN(n_8_0_88));
   INV_X1 i_8_0_102 (.A(n_112), .ZN(n_8_0_89));
   INV_X1 i_8_0_135 (.A(n_71), .ZN(n_8_0_90));
   INV_X1 i_8_0_136 (.A(n_109), .ZN(n_8_0_91));
   INV_X1 i_8_0_137 (.A(n_70), .ZN(n_8_0_92));
   INV_X1 i_8_0_138 (.A(n_107), .ZN(n_8_0_93));
   INV_X1 i_8_0_169 (.A(n_106), .ZN(n_8_0_94));
   INV_X1 i_8_0_170 (.A(n_69), .ZN(n_8_0_95));
   INV_X1 i_8_0_172 (.A(in1[0]), .ZN(n_8_0_96));
   INV_X1 i_8_0_203 (.A(in2[0]), .ZN(n_8_0_97));
   NOR2_X1 i_8_0_204 (.A1(n_8_0_84), .A2(n_8_0_97), .ZN(n_8_25));
   NOR2_X1 i_8_0_237 (.A1(n_8_0_82), .A2(n_8_0_97), .ZN(n_8_27));
   NOR2_X1 i_8_0_238 (.A1(n_8_0_81), .A2(n_8_0_97), .ZN(n_8_28));
   NOR2_X1 i_8_0_239 (.A1(n_8_0_78), .A2(n_8_0_96), .ZN(n_8_65));
   NOR2_X1 i_8_0_240 (.A1(n_8_0_77), .A2(n_8_0_96), .ZN(n_8_98));
   NOR2_X1 i_8_0_271 (.A1(n_8_0_77), .A2(n_8_0_95), .ZN(n_8_99));
   NOR2_X1 i_8_0_273 (.A1(n_8_0_77), .A2(n_8_0_94), .ZN(n_8_100));
   NOR2_X1 i_8_0_274 (.A1(n_8_0_76), .A2(n_8_0_96), .ZN(n_8_131));
   NOR2_X1 i_8_0_275 (.A1(n_8_0_76), .A2(n_8_0_94), .ZN(n_8_133));
   NOR2_X1 i_8_0_276 (.A1(n_8_0_75), .A2(n_8_0_96), .ZN(n_8_164));
   NOR2_X1 i_8_0_278 (.A1(n_8_0_74), .A2(n_8_0_96), .ZN(n_8_197));
   NOR2_X1 i_8_0_280 (.A1(n_8_0_74), .A2(n_8_0_95), .ZN(n_8_198));
   NOR2_X1 i_8_0_282 (.A1(n_8_0_74), .A2(n_8_0_94), .ZN(n_8_199));
   NOR2_X1 i_8_0_283 (.A1(n_8_0_73), .A2(n_8_0_95), .ZN(n_8_231));
   NOR2_X1 i_8_0_284 (.A1(n_8_0_73), .A2(n_8_0_94), .ZN(n_8_232));
   NOR2_X1 i_8_0_815 (.A1(n_8_0_73), .A2(n_8_0_93), .ZN(n_8_233));
   NOR2_X1 i_8_0_845 (.A1(n_8_0_73), .A2(n_8_0_92), .ZN(n_8_234));
   NOR2_X1 i_8_0_849 (.A1(n_8_0_73), .A2(n_8_0_91), .ZN(n_8_236));
   NOR2_X1 i_8_0_878 (.A1(n_8_0_73), .A2(n_8_0_90), .ZN(n_8_238));
   NOR2_X1 i_8_0_880 (.A1(n_8_0_73), .A2(n_8_0_89), .ZN(n_8_240));
   NOR2_X1 i_8_0_883 (.A1(n_8_0_73), .A2(n_8_0_88), .ZN(n_8_241));
   NOR2_X1 i_8_0_913 (.A1(n_8_0_73), .A2(n_8_0_87), .ZN(n_8_242));
   NOR2_X1 i_8_0_915 (.A1(n_8_0_81), .A2(n_8_0_72), .ZN(n_8_505));
   NOR2_X1 i_8_0_917 (.A1(n_8_0_82), .A2(n_8_0_71), .ZN(n_8_448));
   NOR2_X1 i_8_0_947 (.A1(n_8_0_80), .A2(n_8_0_71), .ZN(n_8_450));
   NOR2_X1 i_8_0_948 (.A1(n_8_0_81), .A2(n_8_0_70), .ZN(n_8_460));
   NOR2_X1 i_8_0_950 (.A1(n_8_0_79), .A2(n_8_0_70), .ZN(n_8_462));
   NOR2_X1 i_8_0_951 (.A1(n_8_0_81), .A2(n_8_0_69), .ZN(n_8_527));
   NOR2_X1 i_8_0_983 (.A1(n_8_0_80), .A2(n_8_0_69), .ZN(n_8_528));
   NOR2_X1 i_8_0_984 (.A1(n_8_0_98), .A2(n_8_0_69), .ZN(n_8_530));
   NOR2_X1 i_8_0_985 (.A1(n_8_0_79), .A2(n_8_0_68), .ZN(n_8_627));
   NOR2_X1 i_8_0_1010 (.A1(n_8_0_98), .A2(n_8_0_68), .ZN(n_8_628));
   NOR2_X1 i_8_0_1015 (.A1(n_8_0_86), .A2(n_8_0_99), .ZN(n_8_686));
   NOR2_X1 i_8_0_1018 (.A1(n_8_0_81), .A2(n_8_0_99), .ZN(n_8_724));
   NOR2_X1 i_8_0_1019 (.A1(n_8_0_85), .A2(n_8_0_67), .ZN(n_8_786));
   NOR2_X1 i_8_0_1045 (.A1(n_8_0_81), .A2(n_8_0_67), .ZN(n_8_823));
   NOR2_X1 i_8_0_1049 (.A1(n_8_0_84), .A2(n_8_0_66), .ZN(n_8_887));
   NOR2_X1 i_8_0_1053 (.A1(n_8_0_82), .A2(n_8_0_66), .ZN(n_8_921));
   NOR2_X1 i_8_0_1080 (.A1(n_8_0_83), .A2(n_8_0_65), .ZN(n_8_1019));
   NOR2_X1 i_8_0_1082 (.A1(n_8_0_81), .A2(n_8_0_65), .ZN(n_8_1021));
   BUF_X1 i_8_0_1087 (.A(n_8_0_65), .Z(n_8_0_64));
   BUF_X1 i_8_0_1115 (.A(n_8_0_66), .Z(n_8_0_63));
   BUF_X1 i_8_0_1117 (.A(n_8_0_67), .Z(n_8_0_62));
   BUF_X1 i_8_0_1121 (.A(n_8_0_99), .Z(n_8_0_61));
   BUF_X1 i_8_0_1122 (.A(n_8_0_68), .Z(n_8_0_60));
   BUF_X1 i_8_0_1123 (.A(n_8_0_69), .Z(n_8_0_59));
   BUF_X1 i_8_0_1124 (.A(n_8_0_70), .Z(n_8_0_58));
   BUF_X1 i_8_0_1125 (.A(n_8_0_71), .Z(n_8_0_57));
   BUF_X1 i_8_0_1126 (.A(n_8_0_72), .Z(n_8_0_56));
   BUF_X1 i_8_0_1127 (.A(n_8_0_73), .Z(n_8_0_40));
   BUF_X1 i_8_0_1128 (.A(n_8_0_74), .Z(n_8_0_39));
   BUF_X1 i_8_0_1129 (.A(n_8_0_75), .Z(n_8_0_38));
   BUF_X1 i_8_0_1130 (.A(n_8_0_76), .Z(n_8_0_37));
   BUF_X1 i_8_0_1131 (.A(n_8_0_77), .Z(n_8_0_36));
   BUF_X1 i_8_0_1132 (.A(n_8_0_78), .Z(n_8_0_35));
   BUF_X1 i_8_0_1133 (.A(n_8_0_98), .Z(n_8_0_33));
   BUF_X1 i_8_0_1134 (.A(n_8_0_79), .Z(n_8_0_32));
   BUF_X1 i_8_0_1135 (.A(n_8_0_80), .Z(n_8_0_31));
   BUF_X1 i_8_0_1136 (.A(n_8_0_81), .Z(n_8_0_30));
   BUF_X1 i_8_0_1137 (.A(n_8_0_82), .Z(n_8_0_29));
   BUF_X1 i_8_0_1138 (.A(n_8_0_83), .Z(n_8_0_28));
   BUF_X1 i_8_0_1139 (.A(n_8_0_84), .Z(n_8_0_27));
   BUF_X1 i_8_0_1140 (.A(n_8_0_85), .Z(n_8_0_26));
   BUF_X1 i_8_0_1141 (.A(n_8_0_86), .Z(n_8_0_25));
   BUF_X1 i_8_0_1142 (.A(n_8_0_87), .Z(n_8_0_13));
   BUF_X1 i_8_0_1143 (.A(n_8_0_88), .Z(n_8_0_12));
   BUF_X1 i_8_0_1144 (.A(n_8_0_89), .Z(n_8_0_11));
   BUF_X1 i_8_0_1145 (.A(n_8_0_90), .Z(n_8_0_9));
   BUF_X1 i_8_0_1146 (.A(n_8_0_91), .Z(n_8_0_7));
   BUF_X1 i_8_0_1147 (.A(n_8_0_92), .Z(n_8_0_5));
   BUF_X1 i_8_0_1148 (.A(n_8_0_93), .Z(n_8_0_4));
   BUF_X1 i_8_0_1149 (.A(n_8_0_94), .Z(n_8_0_3));
   BUF_X1 i_8_0_1150 (.A(n_8_0_95), .Z(n_8_0_2));
   BUF_X1 i_8_0_1151 (.A(n_8_0_96), .Z(n_8_0_1));
   BUF_X1 i_8_0_1152 (.A(n_8_0_97), .Z(n_8_0_0));
   INV_X1 i_8_0_1153 (.A(n_76), .ZN(n_8_0_98));
   INV_X1 i_8_0_1154 (.A(n_86), .ZN(n_8_0_99));
   INV_X1 i_8_0_1155 (.A(n_8_0_100), .ZN(n_8_727));
   NAND2_X1 i_8_0_1156 (.A1(n_76), .A2(n_86), .ZN(n_8_0_100));
   datapath__0_65 i_1_6 (.p_0({n_1_30, n_1_29, n_1_28, n_1_27, n_1_26, n_1_25, 
      n_1_24, n_1_23, n_1_22, n_1_21, n_1_20, n_1_19, n_1_18, n_1_17, n_1_16, 
      n_1_15, n_1_14, n_1_13, n_1_12, n_1_11, n_1_10, n_1_9, n_1_8, n_1_7, n_1_6, 
      n_1_5, n_1_4, n_1_3, n_1_2, n_1_1, n_1_0, uc_994}), .in2(in2));
   datapath i_1_1 (.p_0({n_1_61, n_1_60, n_1_59, n_1_58, n_1_57, n_1_56, n_1_55, 
      n_1_54, n_1_53, n_1_52, n_1_51, n_1_50, n_1_49, n_1_48, n_1_47, n_1_46, 
      n_1_45, n_1_44, n_1_43, n_1_42, n_1_41, n_1_40, n_1_39, n_1_38, n_1_37, 
      n_1_36, n_1_35, n_1_34, n_1_33, n_1_32, n_1_31, uc_995}), .in1(in1));
   MUX2_X1 i_1_0_0 (.A(in2[1]), .B(n_1_0), .S(in2[31]), .Z(n_64));
   MUX2_X1 i_1_0_1 (.A(in2[2]), .B(n_1_1), .S(in2[31]), .Z(n_65));
   MUX2_X1 i_1_0_2 (.A(in2[3]), .B(n_1_2), .S(in2[31]), .Z(n_66));
   MUX2_X1 i_1_0_11 (.A(in2[12]), .B(n_1_11), .S(in2[31]), .Z(n_67));
   AND2_X1 i_1_0_30 (.A1(in2[31]), .A2(n_1_30), .ZN(n_68));
   MUX2_X1 i_1_0_31 (.A(in1[1]), .B(n_1_31), .S(in2[31]), .Z(n_69));
   MUX2_X1 i_1_0_34 (.A(in1[4]), .B(n_1_34), .S(in2[31]), .Z(n_70));
   MUX2_X1 i_1_0_38 (.A(in1[8]), .B(n_1_38), .S(in2[31]), .Z(n_71));
   MUX2_X1 i_1_0_53 (.A(in1[23]), .B(n_1_53), .S(in2[31]), .Z(n_72));
   MUX2_X1 i_1_0_55 (.A(in1[25]), .B(n_1_55), .S(in2[31]), .Z(n_73));
   MUX2_X1 i_1_0_58 (.A(in1[28]), .B(n_1_58), .S(in2[31]), .Z(n_74));
   MUX2_X1 i_1_0_60 (.A(in1[30]), .B(n_1_60), .S(in2[31]), .Z(n_75));
   OAI21_X1 i_1_0_61 (.A(n_1_0_0), .B1(n_1_0_1), .B2(in1[31]), .ZN(n_76));
   INV_X1 i_1_0_62 (.A(n_77), .ZN(n_1_0_0));
   MUX2_X1 i_1_0_63 (.A(in1[31]), .B(n_1_61), .S(in2[31]), .Z(n_77));
   INV_X1 i_1_0_64 (.A(in2[31]), .ZN(n_1_0_1));
   OR2_X1 i_1_0_3 (.A1(in2[31]), .A2(in2[28]), .ZN(n_1_0_2));
   OR2_X1 i_1_0_4 (.A1(in2[31]), .A2(in2[29]), .ZN(n_1_0_3));
   OR2_X1 i_1_0_5 (.A1(in2[31]), .A2(in2[30]), .ZN(n_1_0_4));
   OAI21_X1 i_1_0_6 (.A(n_1_0_5), .B1(n_1_0_6), .B2(in2[31]), .ZN(n_78));
   NAND2_X1 i_1_0_7 (.A1(in2[31]), .A2(n_1_22), .ZN(n_1_0_5));
   INV_X1 i_1_0_8 (.A(in2[23]), .ZN(n_1_0_6));
   INV_X1 i_1_0_9 (.A(n_1_0_7), .ZN(n_79));
   OAI21_X1 i_1_0_10 (.A(n_1_0_2), .B1(n_1_0_10), .B2(n_1_27), .ZN(n_1_0_7));
   INV_X1 i_1_0_12 (.A(n_1_0_8), .ZN(n_80));
   OAI21_X1 i_1_0_13 (.A(n_1_0_3), .B1(n_1_0_10), .B2(n_1_28), .ZN(n_1_0_8));
   INV_X1 i_1_0_14 (.A(n_1_0_9), .ZN(n_81));
   OAI21_X1 i_1_0_15 (.A(n_1_0_4), .B1(n_1_0_10), .B2(n_1_29), .ZN(n_1_0_9));
   INV_X1 i_1_0_16 (.A(in2[31]), .ZN(n_1_0_10));
   OAI21_X1 i_1_0_17 (.A(n_1_0_11), .B1(n_1_0_12), .B2(in2[31]), .ZN(n_82));
   NAND2_X1 i_1_0_18 (.A1(in2[31]), .A2(n_1_48), .ZN(n_1_0_11));
   INV_X1 i_1_0_19 (.A(in1[18]), .ZN(n_1_0_12));
   OAI21_X1 i_1_0_20 (.A(n_1_0_13), .B1(n_1_0_14), .B2(in2[31]), .ZN(n_83));
   NAND2_X1 i_1_0_21 (.A1(in2[31]), .A2(n_1_51), .ZN(n_1_0_13));
   INV_X1 i_1_0_22 (.A(in1[21]), .ZN(n_1_0_14));
   OAI21_X1 i_1_0_23 (.A(n_1_0_15), .B1(n_1_0_16), .B2(in2[31]), .ZN(n_84));
   NAND2_X1 i_1_0_24 (.A1(in2[31]), .A2(n_1_54), .ZN(n_1_0_15));
   INV_X1 i_1_0_25 (.A(in1[24]), .ZN(n_1_0_16));
   OAI21_X1 i_1_0_26 (.A(n_1_0_17), .B1(n_1_0_18), .B2(in2[31]), .ZN(n_85));
   NAND2_X1 i_1_0_27 (.A1(in2[31]), .A2(n_1_59), .ZN(n_1_0_17));
   INV_X1 i_1_0_28 (.A(in1[29]), .ZN(n_1_0_18));
   NAND2_X1 i_1_0_29 (.A1(n_1_0_19), .A2(n_1_0_20), .ZN(n_86));
   NAND2_X1 i_1_0_32 (.A1(n_1_0_94), .A2(in2[4]), .ZN(n_1_0_19));
   NAND2_X1 i_1_0_33 (.A1(in2[31]), .A2(n_1_3), .ZN(n_1_0_20));
   NAND2_X1 i_1_0_35 (.A1(n_1_0_21), .A2(n_1_0_22), .ZN(n_87));
   NAND2_X1 i_1_0_36 (.A1(n_1_0_94), .A2(in2[5]), .ZN(n_1_0_21));
   NAND2_X1 i_1_0_37 (.A1(in2[31]), .A2(n_1_4), .ZN(n_1_0_22));
   NAND2_X1 i_1_0_39 (.A1(n_1_0_23), .A2(n_1_0_24), .ZN(n_88));
   NAND2_X1 i_1_0_40 (.A1(n_1_0_94), .A2(in2[6]), .ZN(n_1_0_23));
   NAND2_X1 i_1_0_41 (.A1(in2[31]), .A2(n_1_5), .ZN(n_1_0_24));
   NAND2_X1 i_1_0_42 (.A1(n_1_0_25), .A2(n_1_0_26), .ZN(n_89));
   NAND2_X1 i_1_0_43 (.A1(n_1_0_94), .A2(in2[7]), .ZN(n_1_0_25));
   NAND2_X1 i_1_0_44 (.A1(in2[31]), .A2(n_1_6), .ZN(n_1_0_26));
   NAND2_X1 i_1_0_45 (.A1(n_1_0_27), .A2(n_1_0_28), .ZN(n_90));
   NAND2_X1 i_1_0_46 (.A1(n_1_0_94), .A2(in2[8]), .ZN(n_1_0_27));
   NAND2_X1 i_1_0_47 (.A1(in2[31]), .A2(n_1_7), .ZN(n_1_0_28));
   NAND2_X1 i_1_0_48 (.A1(n_1_0_29), .A2(n_1_0_30), .ZN(n_91));
   NAND2_X1 i_1_0_49 (.A1(n_1_0_94), .A2(in2[9]), .ZN(n_1_0_29));
   NAND2_X1 i_1_0_50 (.A1(in2[31]), .A2(n_1_8), .ZN(n_1_0_30));
   NAND2_X1 i_1_0_51 (.A1(n_1_0_31), .A2(n_1_0_32), .ZN(n_92));
   NAND2_X1 i_1_0_52 (.A1(n_1_0_94), .A2(in2[10]), .ZN(n_1_0_31));
   NAND2_X1 i_1_0_54 (.A1(in2[31]), .A2(n_1_9), .ZN(n_1_0_32));
   NAND2_X1 i_1_0_56 (.A1(n_1_0_33), .A2(n_1_0_34), .ZN(n_93));
   NAND2_X1 i_1_0_57 (.A1(n_1_0_94), .A2(in2[13]), .ZN(n_1_0_33));
   NAND2_X1 i_1_0_59 (.A1(in2[31]), .A2(n_1_12), .ZN(n_1_0_34));
   NAND2_X1 i_1_0_65 (.A1(n_1_0_35), .A2(n_1_0_36), .ZN(n_94));
   NAND2_X1 i_1_0_66 (.A1(n_1_0_94), .A2(in2[15]), .ZN(n_1_0_35));
   NAND2_X1 i_1_0_67 (.A1(in2[31]), .A2(n_1_14), .ZN(n_1_0_36));
   NAND2_X1 i_1_0_68 (.A1(n_1_0_37), .A2(n_1_0_38), .ZN(n_95));
   NAND2_X1 i_1_0_69 (.A1(n_1_0_94), .A2(in2[16]), .ZN(n_1_0_37));
   NAND2_X1 i_1_0_70 (.A1(in2[31]), .A2(n_1_15), .ZN(n_1_0_38));
   NAND2_X1 i_1_0_71 (.A1(n_1_0_39), .A2(n_1_0_40), .ZN(n_96));
   NAND2_X1 i_1_0_72 (.A1(n_1_0_94), .A2(in2[17]), .ZN(n_1_0_39));
   NAND2_X1 i_1_0_73 (.A1(in2[31]), .A2(n_1_16), .ZN(n_1_0_40));
   NAND2_X1 i_1_0_74 (.A1(n_1_0_41), .A2(n_1_0_42), .ZN(n_97));
   NAND2_X1 i_1_0_75 (.A1(n_1_0_94), .A2(in2[18]), .ZN(n_1_0_41));
   NAND2_X1 i_1_0_76 (.A1(in2[31]), .A2(n_1_17), .ZN(n_1_0_42));
   NAND2_X1 i_1_0_77 (.A1(n_1_0_43), .A2(n_1_0_44), .ZN(n_98));
   NAND2_X1 i_1_0_78 (.A1(n_1_0_94), .A2(in2[19]), .ZN(n_1_0_43));
   NAND2_X1 i_1_0_79 (.A1(in2[31]), .A2(n_1_18), .ZN(n_1_0_44));
   NAND2_X1 i_1_0_80 (.A1(n_1_0_45), .A2(n_1_0_46), .ZN(n_99));
   NAND2_X1 i_1_0_81 (.A1(n_1_0_94), .A2(in2[20]), .ZN(n_1_0_45));
   NAND2_X1 i_1_0_82 (.A1(in2[31]), .A2(n_1_19), .ZN(n_1_0_46));
   NAND2_X1 i_1_0_83 (.A1(n_1_0_47), .A2(n_1_0_48), .ZN(n_100));
   NAND2_X1 i_1_0_84 (.A1(n_1_0_94), .A2(in2[21]), .ZN(n_1_0_47));
   NAND2_X1 i_1_0_85 (.A1(in2[31]), .A2(n_1_20), .ZN(n_1_0_48));
   NAND2_X1 i_1_0_86 (.A1(n_1_0_49), .A2(n_1_0_50), .ZN(n_101));
   NAND2_X1 i_1_0_87 (.A1(n_1_0_94), .A2(in2[22]), .ZN(n_1_0_49));
   NAND2_X1 i_1_0_88 (.A1(in2[31]), .A2(n_1_21), .ZN(n_1_0_50));
   NAND2_X1 i_1_0_89 (.A1(n_1_0_51), .A2(n_1_0_52), .ZN(n_102));
   NAND2_X1 i_1_0_90 (.A1(n_1_0_94), .A2(in2[24]), .ZN(n_1_0_51));
   NAND2_X1 i_1_0_91 (.A1(in2[31]), .A2(n_1_23), .ZN(n_1_0_52));
   NAND2_X1 i_1_0_92 (.A1(n_1_0_53), .A2(n_1_0_54), .ZN(n_103));
   NAND2_X1 i_1_0_93 (.A1(n_1_0_94), .A2(in2[25]), .ZN(n_1_0_53));
   NAND2_X1 i_1_0_94 (.A1(in2[31]), .A2(n_1_24), .ZN(n_1_0_54));
   NAND2_X1 i_1_0_95 (.A1(n_1_0_55), .A2(n_1_0_56), .ZN(n_104));
   NAND2_X1 i_1_0_96 (.A1(n_1_0_94), .A2(in2[26]), .ZN(n_1_0_55));
   NAND2_X1 i_1_0_97 (.A1(in2[31]), .A2(n_1_25), .ZN(n_1_0_56));
   NAND2_X1 i_1_0_98 (.A1(n_1_0_57), .A2(n_1_0_58), .ZN(n_105));
   NAND2_X1 i_1_0_99 (.A1(n_1_0_94), .A2(in2[27]), .ZN(n_1_0_57));
   NAND2_X1 i_1_0_100 (.A1(in2[31]), .A2(n_1_26), .ZN(n_1_0_58));
   NAND2_X1 i_1_0_101 (.A1(n_1_0_59), .A2(n_1_0_60), .ZN(n_106));
   NAND2_X1 i_1_0_102 (.A1(n_1_0_94), .A2(in1[2]), .ZN(n_1_0_59));
   NAND2_X1 i_1_0_103 (.A1(in2[31]), .A2(n_1_32), .ZN(n_1_0_60));
   NAND2_X1 i_1_0_104 (.A1(n_1_0_61), .A2(n_1_0_62), .ZN(n_107));
   NAND2_X1 i_1_0_105 (.A1(n_1_0_94), .A2(in1[3]), .ZN(n_1_0_61));
   NAND2_X1 i_1_0_106 (.A1(in2[31]), .A2(n_1_33), .ZN(n_1_0_62));
   NAND2_X1 i_1_0_107 (.A1(n_1_0_63), .A2(n_1_0_64), .ZN(n_108));
   NAND2_X1 i_1_0_108 (.A1(n_1_0_94), .A2(in1[5]), .ZN(n_1_0_63));
   NAND2_X1 i_1_0_109 (.A1(in2[31]), .A2(n_1_35), .ZN(n_1_0_64));
   NAND2_X1 i_1_0_110 (.A1(n_1_0_65), .A2(n_1_0_66), .ZN(n_109));
   NAND2_X1 i_1_0_111 (.A1(n_1_0_94), .A2(in1[6]), .ZN(n_1_0_65));
   NAND2_X1 i_1_0_112 (.A1(in2[31]), .A2(n_1_36), .ZN(n_1_0_66));
   NAND2_X1 i_1_0_113 (.A1(n_1_0_67), .A2(n_1_0_68), .ZN(n_110));
   NAND2_X1 i_1_0_114 (.A1(n_1_0_94), .A2(in1[7]), .ZN(n_1_0_67));
   NAND2_X1 i_1_0_115 (.A1(in2[31]), .A2(n_1_37), .ZN(n_1_0_68));
   NAND2_X1 i_1_0_116 (.A1(n_1_0_69), .A2(n_1_0_70), .ZN(n_111));
   NAND2_X1 i_1_0_117 (.A1(n_1_0_94), .A2(in1[9]), .ZN(n_1_0_69));
   NAND2_X1 i_1_0_118 (.A1(in2[31]), .A2(n_1_39), .ZN(n_1_0_70));
   NAND2_X1 i_1_0_119 (.A1(n_1_0_71), .A2(n_1_0_72), .ZN(n_112));
   NAND2_X1 i_1_0_120 (.A1(n_1_0_94), .A2(in1[10]), .ZN(n_1_0_71));
   NAND2_X1 i_1_0_121 (.A1(in2[31]), .A2(n_1_40), .ZN(n_1_0_72));
   NAND2_X1 i_1_0_122 (.A1(n_1_0_73), .A2(n_1_0_74), .ZN(n_113));
   NAND2_X1 i_1_0_123 (.A1(n_1_0_94), .A2(in1[11]), .ZN(n_1_0_73));
   NAND2_X1 i_1_0_124 (.A1(in2[31]), .A2(n_1_41), .ZN(n_1_0_74));
   NAND2_X1 i_1_0_125 (.A1(n_1_0_75), .A2(n_1_0_76), .ZN(n_114));
   NAND2_X1 i_1_0_126 (.A1(n_1_0_94), .A2(in1[12]), .ZN(n_1_0_75));
   NAND2_X1 i_1_0_127 (.A1(in2[31]), .A2(n_1_42), .ZN(n_1_0_76));
   NAND2_X1 i_1_0_128 (.A1(n_1_0_77), .A2(n_1_0_78), .ZN(n_115));
   NAND2_X1 i_1_0_129 (.A1(n_1_0_94), .A2(in1[13]), .ZN(n_1_0_77));
   NAND2_X1 i_1_0_130 (.A1(in2[31]), .A2(n_1_43), .ZN(n_1_0_78));
   NAND2_X1 i_1_0_131 (.A1(n_1_0_79), .A2(n_1_0_80), .ZN(n_116));
   NAND2_X1 i_1_0_132 (.A1(n_1_0_94), .A2(in1[14]), .ZN(n_1_0_79));
   NAND2_X1 i_1_0_133 (.A1(in2[31]), .A2(n_1_44), .ZN(n_1_0_80));
   NAND2_X1 i_1_0_134 (.A1(n_1_0_81), .A2(n_1_0_82), .ZN(n_117));
   NAND2_X1 i_1_0_135 (.A1(n_1_0_94), .A2(in1[16]), .ZN(n_1_0_81));
   NAND2_X1 i_1_0_136 (.A1(in2[31]), .A2(n_1_46), .ZN(n_1_0_82));
   NAND2_X1 i_1_0_137 (.A1(n_1_0_83), .A2(n_1_0_84), .ZN(n_118));
   NAND2_X1 i_1_0_138 (.A1(n_1_0_94), .A2(in1[17]), .ZN(n_1_0_83));
   NAND2_X1 i_1_0_139 (.A1(in2[31]), .A2(n_1_47), .ZN(n_1_0_84));
   NAND2_X1 i_1_0_140 (.A1(n_1_0_85), .A2(n_1_0_86), .ZN(n_119));
   NAND2_X1 i_1_0_141 (.A1(n_1_0_94), .A2(in1[19]), .ZN(n_1_0_85));
   NAND2_X1 i_1_0_142 (.A1(in2[31]), .A2(n_1_49), .ZN(n_1_0_86));
   NAND2_X1 i_1_0_143 (.A1(n_1_0_87), .A2(n_1_0_88), .ZN(n_120));
   NAND2_X1 i_1_0_144 (.A1(n_1_0_94), .A2(in1[20]), .ZN(n_1_0_87));
   NAND2_X1 i_1_0_145 (.A1(in2[31]), .A2(n_1_50), .ZN(n_1_0_88));
   NAND2_X1 i_1_0_146 (.A1(n_1_0_89), .A2(n_1_0_90), .ZN(n_121));
   NAND2_X1 i_1_0_147 (.A1(n_1_0_94), .A2(in1[22]), .ZN(n_1_0_89));
   NAND2_X1 i_1_0_148 (.A1(in2[31]), .A2(n_1_52), .ZN(n_1_0_90));
   NAND2_X1 i_1_0_149 (.A1(n_1_0_91), .A2(n_1_0_92), .ZN(n_122));
   NAND2_X1 i_1_0_150 (.A1(n_1_0_94), .A2(in1[26]), .ZN(n_1_0_91));
   NAND2_X1 i_1_0_151 (.A1(in2[31]), .A2(n_1_56), .ZN(n_1_0_92));
   NAND2_X1 i_1_0_152 (.A1(n_1_0_93), .A2(n_1_0_95), .ZN(n_123));
   NAND2_X1 i_1_0_153 (.A1(n_1_0_94), .A2(in1[27]), .ZN(n_1_0_93));
   INV_X1 i_1_0_154 (.A(in2[31]), .ZN(n_1_0_94));
   NAND2_X1 i_1_0_155 (.A1(in2[31]), .A2(n_1_57), .ZN(n_1_0_95));
   NAND2_X1 i_1_0_156 (.A1(n_1_0_96), .A2(n_1_0_97), .ZN(n_124));
   NAND2_X1 i_1_0_157 (.A1(n_1_10), .A2(in2[31]), .ZN(n_1_0_96));
   NAND2_X1 i_1_0_158 (.A1(n_1_0_94), .A2(in2[11]), .ZN(n_1_0_97));
   NAND2_X1 i_1_0_159 (.A1(n_1_0_98), .A2(n_1_0_99), .ZN(n_125));
   NAND2_X1 i_1_0_160 (.A1(n_1_13), .A2(in2[31]), .ZN(n_1_0_98));
   NAND2_X1 i_1_0_161 (.A1(n_1_0_94), .A2(in2[14]), .ZN(n_1_0_99));
   NAND2_X1 i_1_0_162 (.A1(n_1_0_100), .A2(n_1_0_101), .ZN(n_126));
   NAND2_X1 i_1_0_163 (.A1(n_1_45), .A2(in2[31]), .ZN(n_1_0_100));
   NAND2_X1 i_1_0_164 (.A1(n_1_0_94), .A2(in1[15]), .ZN(n_1_0_101));
   DFF_X1 \out_reg[0]  (.D(n_63), .CK(clk), .Q(out[0]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_0), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_1), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_2), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_3), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_4), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_5), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_6), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_7), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_8), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_9), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_10), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_11), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_12), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_13), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_14), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_15), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_16), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_17), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_18), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_19), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_20), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_21), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_22), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_23), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_24), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_25), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_26), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_27), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_28), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_29), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[31]  (.D(n_30), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[32]  (.D(n_31), .CK(clk), .Q(out[32]), .QN());
   DFF_X1 \out_reg[33]  (.D(n_32), .CK(clk), .Q(out[33]), .QN());
   DFF_X1 \out_reg[34]  (.D(n_33), .CK(clk), .Q(out[34]), .QN());
   DFF_X1 \out_reg[35]  (.D(n_34), .CK(clk), .Q(out[35]), .QN());
   DFF_X1 \out_reg[36]  (.D(n_35), .CK(clk), .Q(out[36]), .QN());
   DFF_X1 \out_reg[37]  (.D(n_36), .CK(clk), .Q(out[37]), .QN());
   DFF_X1 \out_reg[38]  (.D(n_37), .CK(clk), .Q(out[38]), .QN());
   DFF_X1 \out_reg[39]  (.D(n_38), .CK(clk), .Q(out[39]), .QN());
   DFF_X1 \out_reg[40]  (.D(n_39), .CK(clk), .Q(out[40]), .QN());
   DFF_X1 \out_reg[41]  (.D(n_40), .CK(clk), .Q(out[41]), .QN());
   DFF_X1 \out_reg[42]  (.D(n_41), .CK(clk), .Q(out[42]), .QN());
   DFF_X1 \out_reg[43]  (.D(n_42), .CK(clk), .Q(out[43]), .QN());
   DFF_X1 \out_reg[44]  (.D(n_43), .CK(clk), .Q(out[44]), .QN());
   DFF_X1 \out_reg[45]  (.D(n_44), .CK(clk), .Q(out[45]), .QN());
   DFF_X1 \out_reg[46]  (.D(n_45), .CK(clk), .Q(out[46]), .QN());
   DFF_X1 \out_reg[47]  (.D(n_46), .CK(clk), .Q(out[47]), .QN());
   DFF_X1 \out_reg[48]  (.D(n_47), .CK(clk), .Q(out[48]), .QN());
   DFF_X1 \out_reg[49]  (.D(n_48), .CK(clk), .Q(out[49]), .QN());
   DFF_X1 \out_reg[50]  (.D(n_49), .CK(clk), .Q(out[50]), .QN());
   DFF_X1 \out_reg[51]  (.D(n_50), .CK(clk), .Q(out[51]), .QN());
   DFF_X1 \out_reg[52]  (.D(n_51), .CK(clk), .Q(out[52]), .QN());
   DFF_X1 \out_reg[53]  (.D(n_52), .CK(clk), .Q(out[53]), .QN());
   DFF_X1 \out_reg[54]  (.D(n_53), .CK(clk), .Q(out[54]), .QN());
   DFF_X1 \out_reg[55]  (.D(n_54), .CK(clk), .Q(out[55]), .QN());
   DFF_X1 \out_reg[56]  (.D(n_55), .CK(clk), .Q(out[56]), .QN());
   DFF_X1 \out_reg[57]  (.D(n_56), .CK(clk), .Q(out[57]), .QN());
   DFF_X1 \out_reg[58]  (.D(n_57), .CK(clk), .Q(out[58]), .QN());
   DFF_X1 \out_reg[59]  (.D(n_58), .CK(clk), .Q(out[59]), .QN());
   DFF_X1 \out_reg[60]  (.D(n_59), .CK(clk), .Q(out[60]), .QN());
   DFF_X1 \out_reg[61]  (.D(n_60), .CK(clk), .Q(out[61]), .QN());
   DFF_X1 \out_reg[62]  (.D(n_61), .CK(clk), .Q(out[62]), .QN());
   DFF_X1 \out_reg[63]  (.D(n_62), .CK(clk), .Q(out[63]), .QN());
endmodule

module Register__parameterized0(in, clk, out);
   input [63:0]in;
   input clk;
   output [63:0]out;

   DFF_X1 \out_reg[63]  (.D(in[63]), .CK(clk), .Q(out[63]), .QN());
   DFF_X1 \out_reg[62]  (.D(in[62]), .CK(clk), .Q(out[62]), .QN());
   DFF_X1 \out_reg[61]  (.D(in[61]), .CK(clk), .Q(out[61]), .QN());
   DFF_X1 \out_reg[60]  (.D(in[60]), .CK(clk), .Q(out[60]), .QN());
   DFF_X1 \out_reg[59]  (.D(in[59]), .CK(clk), .Q(out[59]), .QN());
   DFF_X1 \out_reg[58]  (.D(in[58]), .CK(clk), .Q(out[58]), .QN());
   DFF_X1 \out_reg[57]  (.D(in[57]), .CK(clk), .Q(out[57]), .QN());
   DFF_X1 \out_reg[56]  (.D(in[56]), .CK(clk), .Q(out[56]), .QN());
   DFF_X1 \out_reg[55]  (.D(in[55]), .CK(clk), .Q(out[55]), .QN());
   DFF_X1 \out_reg[54]  (.D(in[54]), .CK(clk), .Q(out[54]), .QN());
   DFF_X1 \out_reg[53]  (.D(in[53]), .CK(clk), .Q(out[53]), .QN());
   DFF_X1 \out_reg[52]  (.D(in[52]), .CK(clk), .Q(out[52]), .QN());
   DFF_X1 \out_reg[51]  (.D(in[51]), .CK(clk), .Q(out[51]), .QN());
   DFF_X1 \out_reg[50]  (.D(in[50]), .CK(clk), .Q(out[50]), .QN());
   DFF_X1 \out_reg[49]  (.D(in[49]), .CK(clk), .Q(out[49]), .QN());
   DFF_X1 \out_reg[48]  (.D(in[48]), .CK(clk), .Q(out[48]), .QN());
   DFF_X1 \out_reg[47]  (.D(in[47]), .CK(clk), .Q(out[47]), .QN());
   DFF_X1 \out_reg[46]  (.D(in[46]), .CK(clk), .Q(out[46]), .QN());
   DFF_X1 \out_reg[45]  (.D(in[45]), .CK(clk), .Q(out[45]), .QN());
   DFF_X1 \out_reg[44]  (.D(in[44]), .CK(clk), .Q(out[44]), .QN());
   DFF_X1 \out_reg[43]  (.D(in[43]), .CK(clk), .Q(out[43]), .QN());
   DFF_X1 \out_reg[42]  (.D(in[42]), .CK(clk), .Q(out[42]), .QN());
   DFF_X1 \out_reg[41]  (.D(in[41]), .CK(clk), .Q(out[41]), .QN());
   DFF_X1 \out_reg[40]  (.D(in[40]), .CK(clk), .Q(out[40]), .QN());
   DFF_X1 \out_reg[39]  (.D(in[39]), .CK(clk), .Q(out[39]), .QN());
   DFF_X1 \out_reg[38]  (.D(in[38]), .CK(clk), .Q(out[38]), .QN());
   DFF_X1 \out_reg[37]  (.D(in[37]), .CK(clk), .Q(out[37]), .QN());
   DFF_X1 \out_reg[36]  (.D(in[36]), .CK(clk), .Q(out[36]), .QN());
   DFF_X1 \out_reg[35]  (.D(in[35]), .CK(clk), .Q(out[35]), .QN());
   DFF_X1 \out_reg[34]  (.D(in[34]), .CK(clk), .Q(out[34]), .QN());
   DFF_X1 \out_reg[33]  (.D(in[33]), .CK(clk), .Q(out[33]), .QN());
   DFF_X1 \out_reg[32]  (.D(in[32]), .CK(clk), .Q(out[32]), .QN());
   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module Register__4_0(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module Register(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module SequentialMultiplierIntegerated(in1, in2, clk, out, ovflag);
   input [31:0]in1;
   input [31:0]in2;
   input clk;
   output [63:0]out;
   output ovflag;

   wire [63:0]result;
   wire [31:0]operand2;
   wire [31:0]operand1;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;

   sequential_multiplier sequential_multiplier_inst (.clk(clk), .rst(), .in1(in1), 
      .in2(in2), .out(result));
   Register__parameterized0 Register_inst3 (.in(result), .clk(clk), .out(out));
   Register__4_0 Register_inst2 (.in(in2), .clk(clk), .out(operand2));
   Register Register_inst1 (.in(in1), .clk(clk), .out(operand1));
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(ovflag));
   OAI221_X1 i_0_0_1 (.A(n_0_0_11), .B1(n_0_0_6), .B2(n_0_0_1), .C1(n_0_0_18), 
      .C2(n_0_0_13), .ZN(n_0_0_0));
   NAND4_X1 i_0_0_2 (.A1(n_0_0_5), .A2(n_0_0_4), .A3(n_0_0_3), .A4(n_0_0_2), 
      .ZN(n_0_0_1));
   NOR4_X1 i_0_0_3 (.A1(operand1[18]), .A2(operand1[17]), .A3(operand1[23]), 
      .A4(operand1[20]), .ZN(n_0_0_2));
   NOR4_X1 i_0_0_4 (.A1(operand1[27]), .A2(operand1[24]), .A3(operand1[30]), 
      .A4(operand1[29]), .ZN(n_0_0_3));
   NOR4_X1 i_0_0_5 (.A1(operand1[6]), .A2(operand1[5]), .A3(operand1[3]), 
      .A4(operand1[0]), .ZN(n_0_0_4));
   NOR4_X1 i_0_0_6 (.A1(operand1[10]), .A2(operand1[9]), .A3(operand1[15]), 
      .A4(operand1[12]), .ZN(n_0_0_5));
   NAND4_X1 i_0_0_7 (.A1(n_0_0_10), .A2(n_0_0_9), .A3(n_0_0_8), .A4(n_0_0_7), 
      .ZN(n_0_0_6));
   NOR4_X1 i_0_0_8 (.A1(operand1[19]), .A2(operand1[16]), .A3(operand1[22]), 
      .A4(operand1[21]), .ZN(n_0_0_7));
   NOR4_X1 i_0_0_9 (.A1(operand1[26]), .A2(operand1[25]), .A3(operand1[31]), 
      .A4(operand1[28]), .ZN(n_0_0_8));
   NOR4_X1 i_0_0_10 (.A1(operand1[2]), .A2(operand1[1]), .A3(operand1[7]), 
      .A4(operand1[4]), .ZN(n_0_0_9));
   NOR4_X1 i_0_0_11 (.A1(operand1[11]), .A2(operand1[8]), .A3(operand1[14]), 
      .A4(operand1[13]), .ZN(n_0_0_10));
   XOR2_X1 i_0_0_12 (.A(out[63]), .B(n_0_0_12), .Z(n_0_0_11));
   XOR2_X1 i_0_0_13 (.A(operand2[31]), .B(operand1[31]), .Z(n_0_0_12));
   NAND4_X1 i_0_0_14 (.A1(n_0_0_17), .A2(n_0_0_16), .A3(n_0_0_15), .A4(n_0_0_14), 
      .ZN(n_0_0_13));
   NOR4_X1 i_0_0_15 (.A1(operand2[7]), .A2(operand2[6]), .A3(operand2[5]), 
      .A4(operand2[4]), .ZN(n_0_0_14));
   NOR4_X1 i_0_0_16 (.A1(operand2[3]), .A2(operand2[2]), .A3(operand2[1]), 
      .A4(operand2[0]), .ZN(n_0_0_15));
   NOR4_X1 i_0_0_17 (.A1(operand2[15]), .A2(operand2[14]), .A3(operand2[13]), 
      .A4(operand2[12]), .ZN(n_0_0_16));
   NOR4_X1 i_0_0_18 (.A1(operand2[11]), .A2(operand2[10]), .A3(operand2[9]), 
      .A4(operand2[8]), .ZN(n_0_0_17));
   NAND4_X1 i_0_0_19 (.A1(n_0_0_22), .A2(n_0_0_21), .A3(n_0_0_20), .A4(n_0_0_19), 
      .ZN(n_0_0_18));
   NOR4_X1 i_0_0_20 (.A1(operand2[25]), .A2(operand2[24]), .A3(operand2[27]), 
      .A4(operand2[26]), .ZN(n_0_0_19));
   NOR4_X1 i_0_0_21 (.A1(operand2[29]), .A2(operand2[28]), .A3(operand2[31]), 
      .A4(operand2[30]), .ZN(n_0_0_20));
   NOR4_X1 i_0_0_22 (.A1(operand2[21]), .A2(operand2[20]), .A3(operand2[23]), 
      .A4(operand2[22]), .ZN(n_0_0_21));
   NOR4_X1 i_0_0_23 (.A1(operand2[17]), .A2(operand2[16]), .A3(operand2[19]), 
      .A4(operand2[18]), .ZN(n_0_0_22));
endmodule
