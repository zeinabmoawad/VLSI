/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Nov  5 17:54:15 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3828786562 */

module datapath(in2, in1, p_0);
   input [7:0]in2;
   input [7:0]in1;
   output [8:0]p_0;

   HA_X1 i_0 (.A(in2[0]), .B(in1[0]), .CO(n_0), .S(p_0[0]));
   FA_X1 i_1 (.A(in2[1]), .B(in1[1]), .CI(n_0), .CO(n_1), .S(p_0[1]));
   FA_X1 i_2 (.A(in2[2]), .B(in1[2]), .CI(n_1), .CO(n_2), .S(p_0[2]));
   FA_X1 i_3 (.A(in2[3]), .B(in1[3]), .CI(n_2), .CO(n_3), .S(p_0[3]));
   FA_X1 i_4 (.A(in2[4]), .B(in1[4]), .CI(n_3), .CO(n_4), .S(p_0[4]));
   FA_X1 i_5 (.A(in2[5]), .B(in1[5]), .CI(n_4), .CO(n_5), .S(p_0[5]));
   FA_X1 i_6 (.A(in2[6]), .B(in1[6]), .CI(n_5), .CO(n_6), .S(p_0[6]));
   FA_X1 i_7 (.A(in2[7]), .B(in1[7]), .CI(n_6), .CO(p_0[8]), .S(p_0[7]));
endmodule

module VerilogAdder(in1, in2, sum, carry);
   input [7:0]in1;
   input [7:0]in2;
   output [7:0]sum;
   output carry;

   datapath i_0 (.in2(in2), .in1(in1), .p_0({carry, sum[7], sum[6], sum[5], 
      sum[4], sum[3], sum[2], sum[1], sum[0]}));
endmodule

module datapath__0_2(EB2, EB);
   output [7:0]EB2;
   input [7:0]EB;

   XOR2_X1 i_0 (.A(EB[1]), .B(EB[0]), .Z(EB2[1]));
   AND2_X1 i_1 (.A1(n_5), .A2(n_0), .ZN(EB2[2]));
   OAI21_X1 i_2 (.A(EB[2]), .B1(EB[1]), .B2(EB[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(EB[3]), .B(n_5), .Z(EB2[3]));
   XOR2_X1 i_4 (.A(EB[4]), .B(n_4), .Z(EB2[4]));
   XOR2_X1 i_5 (.A(EB[5]), .B(n_3), .Z(EB2[5]));
   XOR2_X1 i_6 (.A(EB[6]), .B(n_2), .Z(EB2[6]));
   XNOR2_X1 i_7 (.A(EB[7]), .B(n_1), .ZN(EB2[7]));
   NOR2_X1 i_8 (.A1(n_2), .A2(EB[6]), .ZN(n_1));
   OR2_X1 i_9 (.A1(n_3), .A2(EB[5]), .ZN(n_2));
   OR2_X1 i_10 (.A1(n_4), .A2(EB[4]), .ZN(n_3));
   OR2_X1 i_11 (.A1(n_5), .A2(EB[3]), .ZN(n_4));
   OR3_X1 i_12 (.A1(EB[2]), .A2(EB[1]), .A3(EB[0]), .ZN(n_5));
endmodule

module subtractor(EA, EB, S2, B2);
   input [7:0]EA;
   input [7:0]EB;
   output [7:0]S2;
   output B2;

   wire B;
   wire [7:0]S;
   wire [7:0]EB2;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   VerilogAdder rc (.in1(EA), .in2({EB2[7], EB2[6], EB2[5], EB2[4], EB2[3], 
      EB2[2], EB2[1], EB[0]}), .sum({S[7], S[6], S[5], S[4], S[3], S[2], S[1], 
      S2[0]}), .carry(B));
   datapath__0_2 i_3 (.EB2({EB2[7], EB2[6], EB2[5], EB2[4], EB2[3], EB2[2], 
      EB2[1], uc_0}), .EB(EB));
   XOR2_X1 i_0_0 (.A(S[1]), .B(n_0_7), .Z(S2[1]));
   XNOR2_X1 i_0_1 (.A(S[2]), .B(n_0_6), .ZN(S2[2]));
   XOR2_X1 i_0_2 (.A(S[3]), .B(n_0_0), .Z(S2[3]));
   OAI21_X1 i_0_3 (.A(n_0_6), .B1(n_0_8), .B2(B), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(S[4]), .B(n_0_4), .Z(S2[4]));
   XNOR2_X1 i_0_5 (.A(S[5]), .B(n_0_3), .ZN(S2[5]));
   XOR2_X1 i_0_6 (.A(S[6]), .B(n_0_2), .Z(S2[6]));
   XNOR2_X1 i_0_7 (.A(S[7]), .B(n_0_1), .ZN(S2[7]));
   AOI21_X1 i_0_8 (.A(n_0_2), .B1(S[6]), .B2(B2), .ZN(n_0_1));
   OAI21_X1 i_0_9 (.A(n_0_3), .B1(n_0_9), .B2(B), .ZN(n_0_2));
   AOI21_X1 i_0_10 (.A(n_0_4), .B1(S[4]), .B2(B2), .ZN(n_0_3));
   NAND2_X1 i_0_11 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   OAI21_X1 i_0_12 (.A(B2), .B1(S[3]), .B2(S[2]), .ZN(n_0_5));
   OAI21_X1 i_0_13 (.A(B2), .B1(S[1]), .B2(S2[0]), .ZN(n_0_6));
   AND2_X1 i_0_14 (.A1(S2[0]), .A2(B2), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(B), .ZN(B2));
   INV_X1 i_0_16 (.A(S[2]), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(S[5]), .ZN(n_0_9));
endmodule

module Multiplixer__parameterized0__0_193(A, B, Sel, Out);
   input [24:0]A;
   input [24:0]B;
   input Sel;
   output [24:0]Out;

   MUX2_X1 i_0_0 (.A(A[0]), .B(B[0]), .S(Sel), .Z(Out[0]));
   MUX2_X1 i_0_1 (.A(A[1]), .B(B[1]), .S(Sel), .Z(Out[1]));
   MUX2_X1 i_0_2 (.A(A[2]), .B(B[2]), .S(Sel), .Z(Out[2]));
   MUX2_X1 i_0_3 (.A(A[3]), .B(B[3]), .S(Sel), .Z(Out[3]));
   MUX2_X1 i_0_4 (.A(A[4]), .B(B[4]), .S(Sel), .Z(Out[4]));
   MUX2_X1 i_0_5 (.A(A[5]), .B(B[5]), .S(Sel), .Z(Out[5]));
   MUX2_X1 i_0_6 (.A(A[6]), .B(B[6]), .S(Sel), .Z(Out[6]));
   MUX2_X1 i_0_7 (.A(A[7]), .B(B[7]), .S(Sel), .Z(Out[7]));
   MUX2_X1 i_0_8 (.A(A[8]), .B(B[8]), .S(Sel), .Z(Out[8]));
   MUX2_X1 i_0_9 (.A(A[9]), .B(B[9]), .S(Sel), .Z(Out[9]));
   MUX2_X1 i_0_10 (.A(A[10]), .B(B[10]), .S(Sel), .Z(Out[10]));
   MUX2_X1 i_0_11 (.A(A[11]), .B(B[11]), .S(Sel), .Z(Out[11]));
   MUX2_X1 i_0_12 (.A(A[12]), .B(B[12]), .S(Sel), .Z(Out[12]));
   MUX2_X1 i_0_13 (.A(A[13]), .B(B[13]), .S(Sel), .Z(Out[13]));
   MUX2_X1 i_0_14 (.A(A[14]), .B(B[14]), .S(Sel), .Z(Out[14]));
   MUX2_X1 i_0_15 (.A(A[15]), .B(B[15]), .S(Sel), .Z(Out[15]));
   MUX2_X1 i_0_16 (.A(A[16]), .B(B[16]), .S(Sel), .Z(Out[16]));
   MUX2_X1 i_0_17 (.A(A[17]), .B(B[17]), .S(Sel), .Z(Out[17]));
   MUX2_X1 i_0_18 (.A(A[18]), .B(B[18]), .S(Sel), .Z(Out[18]));
   MUX2_X1 i_0_19 (.A(A[19]), .B(B[19]), .S(Sel), .Z(Out[19]));
   MUX2_X1 i_0_20 (.A(A[20]), .B(B[20]), .S(Sel), .Z(Out[20]));
   MUX2_X1 i_0_21 (.A(A[21]), .B(B[21]), .S(Sel), .Z(Out[21]));
   MUX2_X1 i_0_22 (.A(A[22]), .B(B[22]), .S(Sel), .Z(Out[22]));
   MUX2_X1 i_0_23 (.A(A[24]), .B(B[24]), .S(Sel), .Z(Out[24]));
endmodule

module Multiplixer__parameterized0(A, B, Sel, Out);
   input [24:0]A;
   input [24:0]B;
   input Sel;
   output [24:0]Out;

   MUX2_X1 i_0_0 (.A(A[0]), .B(B[0]), .S(Sel), .Z(Out[0]));
   MUX2_X1 i_0_1 (.A(A[1]), .B(B[1]), .S(Sel), .Z(Out[1]));
   MUX2_X1 i_0_2 (.A(A[2]), .B(B[2]), .S(Sel), .Z(Out[2]));
   MUX2_X1 i_0_3 (.A(A[3]), .B(B[3]), .S(Sel), .Z(Out[3]));
   MUX2_X1 i_0_4 (.A(A[4]), .B(B[4]), .S(Sel), .Z(Out[4]));
   MUX2_X1 i_0_5 (.A(A[5]), .B(B[5]), .S(Sel), .Z(Out[5]));
   MUX2_X1 i_0_6 (.A(A[6]), .B(B[6]), .S(Sel), .Z(Out[6]));
   MUX2_X1 i_0_7 (.A(A[7]), .B(B[7]), .S(Sel), .Z(Out[7]));
   MUX2_X1 i_0_8 (.A(A[8]), .B(B[8]), .S(Sel), .Z(Out[8]));
   MUX2_X1 i_0_9 (.A(A[9]), .B(B[9]), .S(Sel), .Z(Out[9]));
   MUX2_X1 i_0_10 (.A(A[10]), .B(B[10]), .S(Sel), .Z(Out[10]));
   MUX2_X1 i_0_11 (.A(A[11]), .B(B[11]), .S(Sel), .Z(Out[11]));
   MUX2_X1 i_0_12 (.A(A[12]), .B(B[12]), .S(Sel), .Z(Out[12]));
   MUX2_X1 i_0_13 (.A(A[13]), .B(B[13]), .S(Sel), .Z(Out[13]));
   MUX2_X1 i_0_14 (.A(A[14]), .B(B[14]), .S(Sel), .Z(Out[14]));
   MUX2_X1 i_0_15 (.A(A[15]), .B(B[15]), .S(Sel), .Z(Out[15]));
   MUX2_X1 i_0_16 (.A(A[16]), .B(B[16]), .S(Sel), .Z(Out[16]));
   MUX2_X1 i_0_17 (.A(A[17]), .B(B[17]), .S(Sel), .Z(Out[17]));
   MUX2_X1 i_0_18 (.A(A[18]), .B(B[18]), .S(Sel), .Z(Out[18]));
   MUX2_X1 i_0_19 (.A(A[19]), .B(B[19]), .S(Sel), .Z(Out[19]));
   MUX2_X1 i_0_20 (.A(A[20]), .B(B[20]), .S(Sel), .Z(Out[20]));
   MUX2_X1 i_0_21 (.A(A[21]), .B(B[21]), .S(Sel), .Z(Out[21]));
   MUX2_X1 i_0_22 (.A(A[22]), .B(B[22]), .S(Sel), .Z(Out[22]));
   MUX2_X1 i_0_23 (.A(A[24]), .B(B[24]), .S(Sel), .Z(Out[24]));
endmodule

module FA__0_122(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_118(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_114(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_110(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA4bit__0_123(in1, in2, cin, sum, cout);
   input [3:0]in1;
   input [3:0]in2;
   input cin;
   output [3:0]sum;
   output cout;

   wire [4:0]carries;

   FA__0_122 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(carries[1]));
   FA__0_118 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(
      carries[1]), .sum(sum[1]), .cout(carries[2]));
   FA__0_114 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(
      carries[2]), .sum(sum[2]), .cout(carries[3]));
   FA__0_110 genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(
      carries[3]), .sum(sum[3]), .cout(cout));
endmodule

module FA__0_139(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_135(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_131(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_127(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA4bit__0_140(in1, in2, cin, sum, cout);
   input [3:0]in1;
   input [3:0]in2;
   input cin;
   output [3:0]sum;
   output cout;

   wire [4:0]carries;

   FA__0_139 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(carries[1]));
   FA__0_135 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(
      carries[1]), .sum(sum[1]), .cout(carries[2]));
   FA__0_131 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(
      carries[2]), .sum(sum[2]), .cout(carries[3]));
   FA__0_127 genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(
      carries[3]), .sum(sum[3]), .cout(cout));
endmodule

module FA__0_156(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_152(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_148(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_144(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA4bit__0_157(in1, in2, cin, sum, cout);
   input [3:0]in1;
   input [3:0]in2;
   input cin;
   output [3:0]sum;
   output cout;

   wire [4:0]carries;

   FA__0_156 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(carries[1]));
   FA__0_152 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(
      carries[1]), .sum(sum[1]), .cout(carries[2]));
   FA__0_148 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(
      carries[2]), .sum(sum[2]), .cout(carries[3]));
   FA__0_144 genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(
      carries[3]), .sum(sum[3]), .cout(cout));
endmodule

module FA__0_173(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_169(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_165(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_161(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA4bit__0_174(in1, in2, cin, sum, cout);
   input [3:0]in1;
   input [3:0]in2;
   input cin;
   output [3:0]sum;
   output cout;

   wire [4:0]carries;

   FA__0_173 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(carries[1]));
   FA__0_169 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(
      carries[1]), .sum(sum[1]), .cout(carries[2]));
   FA__0_165 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(
      carries[2]), .sum(sum[2]), .cout(carries[3]));
   FA__0_161 genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(
      carries[3]), .sum(sum[3]), .cout(cout));
endmodule

module FA__0_190(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_186(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_182(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_178(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA4bit__0_191(in1, in2, cin, sum, cout);
   input [3:0]in1;
   input [3:0]in2;
   input cin;
   output [3:0]sum;
   output cout;

   wire [4:0]carries;

   FA__0_190 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(carries[1]));
   FA__0_186 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(
      carries[1]), .sum(sum[1]), .cout(carries[2]));
   FA__0_182 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(
      carries[2]), .sum(sum[2]), .cout(carries[3]));
   FA__0_178 genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(
      carries[3]), .sum(sum[3]), .cout(cout));
endmodule

module FA__0_98(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(sum));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(cout));
endmodule

module FA__0_102(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA__0_106(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module FA(in1, in2, cin, sum, cout);
   input in1;
   input in2;
   input cin;
   output sum;
   output cout;

   wire w0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(w0));
   XOR2_X1 i_0_1 (.A(cin), .B(w0), .Z(sum));
   AOI22_X1 i_0_2 (.A1(w0), .A2(cin), .B1(in1), .B2(in2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module RCA4bit(in1, in2, cin, sum, cout);
   input [3:0]in1;
   input [3:0]in2;
   input cin;
   output [3:0]sum;
   output cout;

   wire [4:0]carries;

   FA__0_98 genblk1_0_full_adder_inst (.in1(in1[0]), .in2(in2[0]), .cin(), 
      .sum(sum[0]), .cout(carries[1]));
   FA__0_102 genblk1_1_full_adder_inst (.in1(in1[1]), .in2(in2[1]), .cin(
      carries[1]), .sum(sum[1]), .cout(carries[2]));
   FA__0_106 genblk1_2_full_adder_inst (.in1(in1[2]), .in2(in2[2]), .cin(
      carries[2]), .sum(sum[2]), .cout(carries[3]));
   FA genblk1_3_full_adder_inst (.in1(in1[3]), .in2(in2[3]), .cin(carries[3]), 
      .sum(sum[3]), .cout(cout));
endmodule

module HalfAdder__0_51(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_48(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_45(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_42(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module CIN__0_52(sin, cin, cprev, sumout, carryout);
   input [3:0]sin;
   input cin;
   input cprev;
   output [3:0]sumout;
   output carryout;

   wire cwire0;
   wire cwire1;
   wire cwire2;
   wire cwire3;

   HalfAdder__0_51 HA0 (.x(cprev), .y(sin[0]), .z(sumout[0]), .cout(cwire0));
   HalfAdder__0_48 HA1 (.x(cwire0), .y(sin[1]), .z(sumout[1]), .cout(cwire1));
   HalfAdder__0_45 HA2 (.x(cwire1), .y(sin[2]), .z(sumout[2]), .cout(cwire2));
   HalfAdder__0_42 HA3 (.x(cwire2), .y(sin[3]), .z(sumout[3]), .cout(cwire3));
   OR2_X1 i_0_0 (.A1(cwire3), .A2(cin), .ZN(carryout));
endmodule

module HalfAdder__0_65(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_62(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_59(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_56(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module CIN__0_66(sin, cin, cprev, sumout, carryout);
   input [3:0]sin;
   input cin;
   input cprev;
   output [3:0]sumout;
   output carryout;

   wire cwire0;
   wire cwire1;
   wire cwire2;
   wire cwire3;

   HalfAdder__0_65 HA0 (.x(cprev), .y(sin[0]), .z(sumout[0]), .cout(cwire0));
   HalfAdder__0_62 HA1 (.x(cwire0), .y(sin[1]), .z(sumout[1]), .cout(cwire1));
   HalfAdder__0_59 HA2 (.x(cwire1), .y(sin[2]), .z(sumout[2]), .cout(cwire2));
   HalfAdder__0_56 HA3 (.x(cwire2), .y(sin[3]), .z(sumout[3]), .cout(cwire3));
   OR2_X1 i_0_0 (.A1(cwire3), .A2(cin), .ZN(carryout));
endmodule

module HalfAdder__0_79(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_76(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_73(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_70(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module CIN__0_80(sin, cin, cprev, sumout, carryout);
   input [3:0]sin;
   input cin;
   input cprev;
   output [3:0]sumout;
   output carryout;

   wire cwire0;
   wire cwire1;
   wire cwire2;
   wire cwire3;

   HalfAdder__0_79 HA0 (.x(cprev), .y(sin[0]), .z(sumout[0]), .cout(cwire0));
   HalfAdder__0_76 HA1 (.x(cwire0), .y(sin[1]), .z(sumout[1]), .cout(cwire1));
   HalfAdder__0_73 HA2 (.x(cwire1), .y(sin[2]), .z(sumout[2]), .cout(cwire2));
   HalfAdder__0_70 HA3 (.x(cwire2), .y(sin[3]), .z(sumout[3]), .cout(cwire3));
   OR2_X1 i_0_0 (.A1(cwire3), .A2(cin), .ZN(carryout));
endmodule

module HalfAdder__0_93(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_90(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_87(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_84(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module CIN__0_94(sin, cin, cprev, sumout, carryout);
   input [3:0]sin;
   input cin;
   input cprev;
   output [3:0]sumout;
   output carryout;

   wire cwire0;
   wire cwire1;
   wire cwire2;
   wire cwire3;

   HalfAdder__0_93 HA0 (.x(cprev), .y(sin[0]), .z(sumout[0]), .cout(cwire0));
   HalfAdder__0_90 HA1 (.x(cwire0), .y(sin[1]), .z(sumout[1]), .cout(cwire1));
   HalfAdder__0_87 HA2 (.x(cwire1), .y(sin[2]), .z(sumout[2]), .cout(cwire2));
   HalfAdder__0_84 HA3 (.x(cwire2), .y(sin[3]), .z(sumout[3]), .cout(cwire3));
   OR2_X1 i_0_0 (.A1(cwire3), .A2(cin), .ZN(carryout));
endmodule

module HalfAdder__0_32(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_35(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder__0_38(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module HalfAdder(x, y, z, cout);
   input x;
   input y;
   output z;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(z));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module CIN(sin, cin, cprev, sumout, carryout);
   input [3:0]sin;
   input cin;
   input cprev;
   output [3:0]sumout;
   output carryout;

   wire cwire0;
   wire cwire1;
   wire cwire2;
   wire cwire3;

   HalfAdder__0_32 HA0 (.x(cprev), .y(sin[0]), .z(sumout[0]), .cout(cwire0));
   HalfAdder__0_35 HA1 (.x(cwire0), .y(sin[1]), .z(sumout[1]), .cout(cwire1));
   HalfAdder__0_38 HA2 (.x(cwire1), .y(sin[2]), .z(sumout[2]), .cout(cwire2));
   HalfAdder HA3 (.x(cwire2), .y(sin[3]), .z(sumout[3]), .cout(cwire3));
   OR2_X1 i_0_0 (.A1(cwire3), .A2(cin), .ZN(carryout));
endmodule

module CIA_24bit(in1, in2, sum, carry);
   input [23:0]in1;
   input [23:0]in2;
   output [23:0]sum;
   output carry;

   wire [5:0]carrywire;
   wire [3:0]sumwire5;
   wire [3:0]sumwire4;
   wire [3:0]sumwire3;
   wire [3:0]sumwire2;
   wire [3:0]sumwire1;

   RCA4bit__0_123 RCA5 (.in1({in1[23], in1[22], in1[21], in1[20]}), .in2({
      in2[23], in2[22], in2[21], in2[20]}), .cin(), .sum(sumwire5), .cout(
      carrywire[5]));
   RCA4bit__0_140 RCA4 (.in1({in1[19], in1[18], in1[17], in1[16]}), .in2({
      in2[19], in2[18], in2[17], in2[16]}), .cin(), .sum(sumwire4), .cout(
      carrywire[4]));
   RCA4bit__0_157 RCA3 (.in1({in1[15], in1[14], in1[13], in1[12]}), .in2({
      in2[15], in2[14], in2[13], in2[12]}), .cin(), .sum(sumwire3), .cout(
      carrywire[3]));
   RCA4bit__0_174 RCA2 (.in1({in1[11], in1[10], in1[9], in1[8]}), .in2({in2[11], 
      in2[10], in2[9], in2[8]}), .cin(), .sum(sumwire2), .cout(carrywire[2]));
   RCA4bit__0_191 RCA1 (.in1({in1[7], in1[6], in1[5], in1[4]}), .in2({in2[7], 
      in2[6], in2[5], in2[4]}), .cin(), .sum(sumwire1), .cout(carrywire[1]));
   RCA4bit RCA0 (.in1({in1[3], in1[2], in1[1], in1[0]}), .in2({in2[3], in2[2], 
      in2[1], in2[0]}), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(
      carrywire[0]));
   CIN__0_52 CIN3_4 (.sin(sumwire4), .cin(carrywire[4]), .cprev(n_1), .sumout({
      sum[19], sum[18], sum[17], sum[16]}), .carryout(n_0));
   CIN__0_66 CIN2_3 (.sin(sumwire3), .cin(carrywire[3]), .cprev(n_2), .sumout({
      sum[15], sum[14], sum[13], sum[12]}), .carryout(n_1));
   CIN__0_80 CIN1_2 (.sin(sumwire2), .cin(carrywire[2]), .cprev(n_3), .sumout({
      sum[11], sum[10], sum[9], sum[8]}), .carryout(n_2));
   CIN__0_94 CIN0_1 (.sin(sumwire1), .cin(carrywire[1]), .cprev(carrywire[0]), 
      .sumout({sum[7], sum[6], sum[5], sum[4]}), .carryout(n_3));
   CIN CIN4_5 (.sin(sumwire5), .cin(carrywire[5]), .cprev(n_0), .sumout({sum[23], 
      sum[22], sum[21], sum[20]}), .carryout(carry));
endmodule

module Multiplixer(A, B, Sel, Out);
   input [7:0]A;
   input [7:0]B;
   input Sel;
   output [7:0]Out;

   MUX2_X1 i_0_0 (.A(A[0]), .B(B[0]), .S(Sel), .Z(Out[0]));
   MUX2_X1 i_0_1 (.A(A[1]), .B(B[1]), .S(Sel), .Z(Out[1]));
   MUX2_X1 i_0_2 (.A(A[2]), .B(B[2]), .S(Sel), .Z(Out[2]));
   MUX2_X1 i_0_3 (.A(A[3]), .B(B[3]), .S(Sel), .Z(Out[3]));
   MUX2_X1 i_0_4 (.A(A[4]), .B(B[4]), .S(Sel), .Z(Out[4]));
   MUX2_X1 i_0_5 (.A(A[5]), .B(B[5]), .S(Sel), .Z(Out[5]));
   MUX2_X1 i_0_6 (.A(A[6]), .B(B[6]), .S(Sel), .Z(Out[6]));
   MUX2_X1 i_0_7 (.A(A[7]), .B(B[7]), .S(Sel), .Z(Out[7]));
endmodule

module LZeros(in, out);
   input [23:0]in;
   output [4:0]out;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_10), .B2(in[23]), .ZN(out[0]));
   OAI21_X1 i_0_1 (.A(n_0_9), .B1(n_0_1), .B2(in[16]), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(in[15]), .A2(n_0_2), .ZN(n_0_1));
   AOI21_X1 i_0_3 (.A(in[14]), .B1(n_0_41), .B2(n_0_3), .ZN(n_0_2));
   OAI21_X1 i_0_4 (.A(n_0_40), .B1(in[11]), .B2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(in[10]), .B1(n_0_39), .B2(n_0_5), .ZN(n_0_4));
   OAI21_X1 i_0_6 (.A(n_0_38), .B1(in[7]), .B2(n_0_6), .ZN(n_0_5));
   AOI21_X1 i_0_7 (.A(in[6]), .B1(n_0_37), .B2(n_0_7), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_36), .B1(in[3]), .B2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(in[2]), .B1(n_0_35), .B2(in[0]), .ZN(n_0_8));
   NOR4_X1 i_0_10 (.A1(in[23]), .A2(in[21]), .A3(in[19]), .A4(in[17]), .ZN(n_0_9));
   NOR2_X1 i_0_11 (.A1(in[22]), .A2(n_0_11), .ZN(n_0_10));
   NOR2_X1 i_0_12 (.A1(in[21]), .A2(n_0_12), .ZN(n_0_11));
   AOI21_X1 i_0_13 (.A(in[20]), .B1(n_0_42), .B2(in[18]), .ZN(n_0_12));
   NOR3_X1 i_0_14 (.A1(in[23]), .A2(in[22]), .A3(n_0_13), .ZN(out[1]));
   NOR3_X1 i_0_15 (.A1(in[21]), .A2(in[20]), .A3(n_0_14), .ZN(n_0_13));
   NOR3_X1 i_0_16 (.A1(in[19]), .A2(in[18]), .A3(n_0_15), .ZN(n_0_14));
   NOR3_X1 i_0_17 (.A1(in[17]), .A2(in[16]), .A3(n_0_16), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(in[15]), .A2(in[14]), .A3(n_0_17), .ZN(n_0_16));
   NOR3_X1 i_0_19 (.A1(in[13]), .A2(in[12]), .A3(n_0_18), .ZN(n_0_17));
   NOR3_X1 i_0_20 (.A1(in[11]), .A2(in[10]), .A3(n_0_19), .ZN(n_0_18));
   NOR3_X1 i_0_21 (.A1(in[9]), .A2(in[8]), .A3(n_0_20), .ZN(n_0_19));
   NOR3_X1 i_0_22 (.A1(in[7]), .A2(in[6]), .A3(n_0_21), .ZN(n_0_20));
   NOR3_X1 i_0_23 (.A1(in[5]), .A2(in[4]), .A3(n_0_22), .ZN(n_0_21));
   NOR3_X1 i_0_24 (.A1(in[3]), .A2(in[2]), .A3(n_0_26), .ZN(n_0_22));
   AOI21_X1 i_0_25 (.A(n_0_33), .B1(n_0_23), .B2(n_0_32), .ZN(out[2]));
   NAND2_X1 i_0_26 (.A1(n_0_24), .A2(n_0_30), .ZN(n_0_23));
   OAI21_X1 i_0_27 (.A(n_0_29), .B1(n_0_27), .B2(n_0_25), .ZN(n_0_24));
   AOI21_X1 i_0_28 (.A(n_0_31), .B1(n_0_30), .B2(n_0_29), .ZN(out[3]));
   AOI211_X1 i_0_29 (.A(n_0_31), .B(n_0_28), .C1(n_0_43), .C2(n_0_25), .ZN(
      out[4]));
   NOR4_X1 i_0_30 (.A1(in[3]), .A2(in[2]), .A3(in[1]), .A4(in[0]), .ZN(n_0_25));
   NOR2_X1 i_0_31 (.A1(in[1]), .A2(in[0]), .ZN(n_0_26));
   OR4_X1 i_0_32 (.A1(in[7]), .A2(in[6]), .A3(in[5]), .A4(in[4]), .ZN(n_0_27));
   NAND2_X1 i_0_33 (.A1(n_0_30), .A2(n_0_29), .ZN(n_0_28));
   NOR4_X1 i_0_34 (.A1(in[11]), .A2(in[10]), .A3(in[9]), .A4(in[8]), .ZN(n_0_29));
   NOR4_X1 i_0_35 (.A1(in[15]), .A2(in[14]), .A3(in[13]), .A4(in[12]), .ZN(
      n_0_30));
   NAND2_X1 i_0_36 (.A1(n_0_34), .A2(n_0_32), .ZN(n_0_31));
   NOR4_X1 i_0_37 (.A1(in[19]), .A2(in[18]), .A3(in[17]), .A4(in[16]), .ZN(
      n_0_32));
   INV_X1 i_0_38 (.A(n_0_34), .ZN(n_0_33));
   NOR4_X1 i_0_39 (.A1(in[23]), .A2(in[22]), .A3(in[21]), .A4(in[20]), .ZN(
      n_0_34));
   INV_X1 i_0_40 (.A(in[1]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(in[4]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(in[5]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(in[8]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(in[9]), .ZN(n_0_39));
   INV_X1 i_0_45 (.A(in[12]), .ZN(n_0_40));
   INV_X1 i_0_46 (.A(in[13]), .ZN(n_0_41));
   INV_X1 i_0_47 (.A(in[19]), .ZN(n_0_42));
   INV_X1 i_0_48 (.A(n_0_27), .ZN(n_0_43));
endmodule

module datapath__0_11(p_0, unNormalizedSum);
   output [23:0]p_0;
   input [23:0]unNormalizedSum;

   XOR2_X1 i_0 (.A(unNormalizedSum[1]), .B(unNormalizedSum[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_21), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(unNormalizedSum[2]), .B1(unNormalizedSum[1]), .B2(
      unNormalizedSum[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(unNormalizedSum[3]), .B(n_21), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(unNormalizedSum[4]), .B(n_20), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(unNormalizedSum[5]), .B(n_19), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_18), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(unNormalizedSum[6]), .B1(n_19), .B2(unNormalizedSum[5]), 
      .ZN(n_1));
   XOR2_X1 i_8 (.A(unNormalizedSum[7]), .B(n_18), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(unNormalizedSum[8]), .B(n_17), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_16), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(unNormalizedSum[9]), .B1(n_17), .B2(unNormalizedSum[8]), 
      .ZN(n_2));
   XOR2_X1 i_12 (.A(unNormalizedSum[10]), .B(n_16), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(unNormalizedSum[11]), .B(n_15), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(unNormalizedSum[12]), .B(n_14), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(unNormalizedSum[13]), .B(n_13), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(unNormalizedSum[14]), .B(n_12), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(unNormalizedSum[15]), .B(n_11), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(unNormalizedSum[16]), .B(n_10), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(unNormalizedSum[17]), .B(n_9), .Z(p_0[17]));
   XOR2_X1 i_20 (.A(unNormalizedSum[18]), .B(n_8), .Z(p_0[18]));
   AND2_X1 i_21 (.A1(n_7), .A2(n_3), .ZN(p_0[19]));
   OAI21_X1 i_22 (.A(unNormalizedSum[19]), .B1(n_8), .B2(unNormalizedSum[18]), 
      .ZN(n_3));
   XOR2_X1 i_23 (.A(unNormalizedSum[20]), .B(n_7), .Z(p_0[20]));
   XNOR2_X1 i_24 (.A(unNormalizedSum[21]), .B(n_6), .ZN(p_0[21]));
   XNOR2_X1 i_25 (.A(unNormalizedSum[22]), .B(n_5), .ZN(p_0[22]));
   XNOR2_X1 i_26 (.A(unNormalizedSum[23]), .B(n_4), .ZN(p_0[23]));
   NOR4_X1 i_27 (.A1(n_7), .A2(unNormalizedSum[20]), .A3(unNormalizedSum[21]), 
      .A4(unNormalizedSum[22]), .ZN(n_4));
   NOR3_X1 i_28 (.A1(n_7), .A2(unNormalizedSum[20]), .A3(unNormalizedSum[21]), 
      .ZN(n_5));
   NOR2_X1 i_29 (.A1(n_7), .A2(unNormalizedSum[20]), .ZN(n_6));
   OR3_X1 i_30 (.A1(n_8), .A2(unNormalizedSum[18]), .A3(unNormalizedSum[19]), 
      .ZN(n_7));
   OR2_X1 i_31 (.A1(n_9), .A2(unNormalizedSum[17]), .ZN(n_8));
   OR2_X1 i_32 (.A1(n_10), .A2(unNormalizedSum[16]), .ZN(n_9));
   NAND2_X1 i_33 (.A1(n_11), .A2(n_23), .ZN(n_10));
   NOR3_X1 i_34 (.A1(n_13), .A2(unNormalizedSum[13]), .A3(unNormalizedSum[14]), 
      .ZN(n_11));
   NOR2_X1 i_35 (.A1(n_13), .A2(unNormalizedSum[13]), .ZN(n_12));
   OR2_X1 i_36 (.A1(n_14), .A2(unNormalizedSum[12]), .ZN(n_13));
   NAND2_X1 i_37 (.A1(n_15), .A2(n_22), .ZN(n_14));
   NOR2_X1 i_38 (.A1(n_16), .A2(unNormalizedSum[10]), .ZN(n_15));
   OR3_X1 i_39 (.A1(n_17), .A2(unNormalizedSum[8]), .A3(unNormalizedSum[9]), 
      .ZN(n_16));
   OR2_X1 i_40 (.A1(n_18), .A2(unNormalizedSum[7]), .ZN(n_17));
   OR3_X1 i_41 (.A1(n_19), .A2(unNormalizedSum[5]), .A3(unNormalizedSum[6]), 
      .ZN(n_18));
   OR2_X1 i_42 (.A1(n_20), .A2(unNormalizedSum[4]), .ZN(n_19));
   OR2_X1 i_43 (.A1(n_21), .A2(unNormalizedSum[3]), .ZN(n_20));
   OR3_X1 i_44 (.A1(unNormalizedSum[2]), .A2(unNormalizedSum[1]), .A3(
      unNormalizedSum[0]), .ZN(n_21));
   INV_X1 i_45 (.A(unNormalizedSum[11]), .ZN(n_22));
   INV_X1 i_46 (.A(unNormalizedSum[15]), .ZN(n_23));
endmodule

module datapath__0_24(p_0, shiftedToAdd);
   output [23:0]p_0;
   input [23:0]shiftedToAdd;

   XOR2_X1 i_0 (.A(shiftedToAdd[1]), .B(shiftedToAdd[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_21), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(shiftedToAdd[2]), .B1(shiftedToAdd[1]), .B2(shiftedToAdd[0]), 
      .ZN(n_0));
   XOR2_X1 i_3 (.A(shiftedToAdd[3]), .B(n_21), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(shiftedToAdd[4]), .B(n_20), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(shiftedToAdd[5]), .B(n_19), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_18), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(shiftedToAdd[6]), .B1(n_19), .B2(shiftedToAdd[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(shiftedToAdd[7]), .B(n_18), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(shiftedToAdd[8]), .B(n_17), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_16), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(shiftedToAdd[9]), .B1(n_17), .B2(shiftedToAdd[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(shiftedToAdd[10]), .B(n_16), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(shiftedToAdd[11]), .B(n_15), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(shiftedToAdd[12]), .B(n_14), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(shiftedToAdd[13]), .B(n_13), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(shiftedToAdd[14]), .B(n_12), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(shiftedToAdd[15]), .B(n_11), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(shiftedToAdd[16]), .B(n_10), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(shiftedToAdd[17]), .B(n_9), .Z(p_0[17]));
   XOR2_X1 i_20 (.A(shiftedToAdd[18]), .B(n_8), .Z(p_0[18]));
   AND2_X1 i_21 (.A1(n_7), .A2(n_3), .ZN(p_0[19]));
   OAI21_X1 i_22 (.A(shiftedToAdd[19]), .B1(n_8), .B2(shiftedToAdd[18]), 
      .ZN(n_3));
   XOR2_X1 i_23 (.A(shiftedToAdd[20]), .B(n_7), .Z(p_0[20]));
   XNOR2_X1 i_24 (.A(shiftedToAdd[21]), .B(n_6), .ZN(p_0[21]));
   XNOR2_X1 i_25 (.A(shiftedToAdd[22]), .B(n_5), .ZN(p_0[22]));
   XNOR2_X1 i_26 (.A(shiftedToAdd[23]), .B(n_4), .ZN(p_0[23]));
   NOR4_X1 i_27 (.A1(n_7), .A2(shiftedToAdd[20]), .A3(shiftedToAdd[21]), 
      .A4(shiftedToAdd[22]), .ZN(n_4));
   NOR3_X1 i_28 (.A1(n_7), .A2(shiftedToAdd[20]), .A3(shiftedToAdd[21]), 
      .ZN(n_5));
   NOR2_X1 i_29 (.A1(n_7), .A2(shiftedToAdd[20]), .ZN(n_6));
   OR3_X1 i_30 (.A1(n_8), .A2(shiftedToAdd[18]), .A3(shiftedToAdd[19]), .ZN(n_7));
   OR2_X1 i_31 (.A1(n_9), .A2(shiftedToAdd[17]), .ZN(n_8));
   OR2_X1 i_32 (.A1(n_10), .A2(shiftedToAdd[16]), .ZN(n_9));
   NAND2_X1 i_33 (.A1(n_11), .A2(n_23), .ZN(n_10));
   NOR3_X1 i_34 (.A1(n_13), .A2(shiftedToAdd[13]), .A3(shiftedToAdd[14]), 
      .ZN(n_11));
   NOR2_X1 i_35 (.A1(n_13), .A2(shiftedToAdd[13]), .ZN(n_12));
   OR2_X1 i_36 (.A1(n_14), .A2(shiftedToAdd[12]), .ZN(n_13));
   NAND2_X1 i_37 (.A1(n_15), .A2(n_22), .ZN(n_14));
   NOR2_X1 i_38 (.A1(n_16), .A2(shiftedToAdd[10]), .ZN(n_15));
   OR3_X1 i_39 (.A1(n_17), .A2(shiftedToAdd[8]), .A3(shiftedToAdd[9]), .ZN(n_16));
   OR2_X1 i_40 (.A1(n_18), .A2(shiftedToAdd[7]), .ZN(n_17));
   OR3_X1 i_41 (.A1(n_19), .A2(shiftedToAdd[5]), .A3(shiftedToAdd[6]), .ZN(n_18));
   OR2_X1 i_42 (.A1(n_20), .A2(shiftedToAdd[4]), .ZN(n_19));
   OR2_X1 i_43 (.A1(n_21), .A2(shiftedToAdd[3]), .ZN(n_20));
   OR3_X1 i_44 (.A1(shiftedToAdd[2]), .A2(shiftedToAdd[1]), .A3(shiftedToAdd[0]), 
      .ZN(n_21));
   INV_X1 i_45 (.A(shiftedToAdd[11]), .ZN(n_22));
   INV_X1 i_46 (.A(shiftedToAdd[15]), .ZN(n_23));
endmodule

module datapath__0_27(p_0, outToAdd);
   output [23:0]p_0;
   input [23:0]outToAdd;

   XOR2_X1 i_0 (.A(outToAdd[1]), .B(outToAdd[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_20), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(outToAdd[2]), .B1(outToAdd[1]), .B2(outToAdd[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(outToAdd[3]), .B(n_20), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(outToAdd[4]), .B(n_19), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(outToAdd[5]), .B(n_18), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_17), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(outToAdd[6]), .B1(n_18), .B2(outToAdd[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(outToAdd[7]), .B(n_17), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(outToAdd[8]), .B(n_16), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_15), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(outToAdd[9]), .B1(n_16), .B2(outToAdd[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(outToAdd[10]), .B(n_15), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(outToAdd[11]), .B(n_14), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(outToAdd[12]), .B(n_13), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(outToAdd[13]), .B(n_12), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(outToAdd[14]), .B(n_11), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(outToAdd[15]), .B(n_10), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(outToAdd[16]), .B(n_9), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(outToAdd[17]), .B(n_8), .Z(p_0[17]));
   XNOR2_X1 i_20 (.A(outToAdd[18]), .B(n_7), .ZN(p_0[18]));
   XNOR2_X1 i_21 (.A(outToAdd[19]), .B(n_6), .ZN(p_0[19]));
   XOR2_X1 i_22 (.A(outToAdd[20]), .B(n_5), .Z(p_0[20]));
   XOR2_X1 i_23 (.A(outToAdd[21]), .B(n_4), .Z(p_0[21]));
   XNOR2_X1 i_24 (.A(outToAdd[22]), .B(n_3), .ZN(p_0[22]));
   NOR3_X1 i_25 (.A1(n_4), .A2(outToAdd[21]), .A3(outToAdd[22]), .ZN(p_0[23]));
   NOR2_X1 i_26 (.A1(n_4), .A2(outToAdd[21]), .ZN(n_3));
   OR2_X1 i_27 (.A1(n_5), .A2(outToAdd[20]), .ZN(n_4));
   NAND2_X1 i_28 (.A1(n_6), .A2(n_23), .ZN(n_5));
   NOR3_X1 i_29 (.A1(n_8), .A2(outToAdd[17]), .A3(outToAdd[18]), .ZN(n_6));
   NOR2_X1 i_30 (.A1(n_8), .A2(outToAdd[17]), .ZN(n_7));
   OR2_X1 i_31 (.A1(n_9), .A2(outToAdd[16]), .ZN(n_8));
   NAND2_X1 i_32 (.A1(n_10), .A2(n_22), .ZN(n_9));
   NOR3_X1 i_33 (.A1(n_12), .A2(outToAdd[13]), .A3(outToAdd[14]), .ZN(n_10));
   NOR2_X1 i_34 (.A1(n_12), .A2(outToAdd[13]), .ZN(n_11));
   OR2_X1 i_35 (.A1(n_13), .A2(outToAdd[12]), .ZN(n_12));
   NAND2_X1 i_36 (.A1(n_14), .A2(n_21), .ZN(n_13));
   NOR2_X1 i_37 (.A1(n_15), .A2(outToAdd[10]), .ZN(n_14));
   OR3_X1 i_38 (.A1(n_16), .A2(outToAdd[8]), .A3(outToAdd[9]), .ZN(n_15));
   OR2_X1 i_39 (.A1(n_17), .A2(outToAdd[7]), .ZN(n_16));
   OR3_X1 i_40 (.A1(n_18), .A2(outToAdd[5]), .A3(outToAdd[6]), .ZN(n_17));
   OR2_X1 i_41 (.A1(n_19), .A2(outToAdd[4]), .ZN(n_18));
   OR2_X1 i_42 (.A1(n_20), .A2(outToAdd[3]), .ZN(n_19));
   OR3_X1 i_43 (.A1(outToAdd[2]), .A2(outToAdd[1]), .A3(outToAdd[0]), .ZN(n_20));
   INV_X1 i_44 (.A(outToAdd[11]), .ZN(n_21));
   INV_X1 i_45 (.A(outToAdd[15]), .ZN(n_22));
   INV_X1 i_46 (.A(outToAdd[19]), .ZN(n_23));
endmodule

module floatingadder(a, b, sum, carry);
   input [31:0]a;
   input [31:0]b;
   output [31:0]sum;
   output carry;

   wire borrow;
   wire [7:0]subsum;
   wire [24:0]outToAdd;
   wire [24:0]outToShift;
   wire carryOfM;
   wire [23:0]unNormalizedSum;
   wire [7:0]ES;
   wire [4:0]shiftleftamount;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_1_14;
   wire n_0_1_0;
   wire n_0_1_15;
   wire n_0_1_1;
   wire n_0_1_16;
   wire n_0_1_2;
   wire n_0_1_17;
   wire n_0_1_3;
   wire n_0_1_18;
   wire n_0_1_4;
   wire n_0_1_19;
   wire n_0_1_5;
   wire n_0_1_20;
   wire n_0_1_6;
   wire n_0_1_21;
   wire n_0_1_7;
   wire n_0_1_22;
   wire n_0_1_8;
   wire n_0_1_23;
   wire n_0_1_9;
   wire n_0_1_24;
   wire n_0_1_10;
   wire n_0_1_25;
   wire n_0_1_11;
   wire n_0_1_26;
   wire n_0_1_12;
   wire n_0_1_27;
   wire n_0_1_13;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_1_32;
   wire [23:0]comB;
   wire [23:0]comA;
   wire n_0_1_33;
   wire n_0_1_34;
   wire n_0_1_35;
   wire n_0_1_36;
   wire n_0_1_37;
   wire n_0_1_38;
   wire n_0_1_39;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_1_42;
   wire n_0_1_43;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_1_46;
   wire n_0_1_47;
   wire n_0_1_48;
   wire n_0_1_49;
   wire n_0_1_50;
   wire n_0_1_51;
   wire n_0_1_52;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_61;
   wire n_0_1_62;
   wire n_0_1_63;
   wire n_0_1_64;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_1_104;
   wire n_0_1_105;
   wire n_0_1_106;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_1_113;
   wire n_0_1_114;
   wire n_0_1_115;
   wire n_0_1_116;
   wire n_0_1_117;
   wire n_0_1_118;
   wire n_0_1_119;
   wire n_0_1_120;
   wire n_0_1_121;
   wire n_0_1_122;
   wire n_0_1_123;
   wire n_0_1_124;
   wire n_0_1_125;
   wire n_0_1_126;
   wire n_0_1_127;
   wire n_0_1_128;
   wire n_0_1_129;
   wire n_0_1_130;
   wire n_0_1_131;
   wire n_0_1_132;
   wire n_0_1_133;
   wire n_0_1_134;
   wire n_0_1_135;
   wire n_0_1_136;
   wire n_0_1_137;
   wire n_0_1_138;
   wire n_0_1_139;
   wire n_0_1_140;
   wire n_0_1_141;
   wire n_0_1_142;
   wire n_0_1_143;
   wire n_0_1_144;
   wire n_0_1_145;
   wire n_0_1_146;
   wire n_0_1_147;
   wire n_0_1_148;
   wire n_0_1_149;
   wire n_0_1_150;
   wire n_0_1_151;
   wire n_0_1_152;
   wire n_0_1_153;
   wire n_0_1_154;
   wire n_0_1_155;
   wire n_0_1_156;
   wire n_0_1_157;
   wire n_0_1_158;
   wire n_0_1_159;
   wire n_0_1_160;
   wire n_0_1_161;
   wire n_0_1_162;
   wire n_0_1_163;
   wire n_0_1_164;
   wire n_0_1_165;
   wire n_0_1_166;
   wire n_0_1_167;
   wire n_0_1_168;
   wire n_0_1_169;
   wire n_0_1_170;
   wire n_0_1_171;
   wire n_0_1_172;
   wire n_0_1_173;
   wire n_0_1_174;
   wire n_0_1_175;
   wire n_0_1_176;
   wire n_0_1_177;
   wire n_0_1_178;
   wire n_0_1_179;
   wire [23:0]unNormalizedSum2;
   wire n_0_1_180;
   wire n_0_1_181;
   wire n_0_1_182;
   wire n_0_1_183;
   wire n_0_1_184;
   wire n_0_1_185;
   wire n_0_1_186;
   wire n_0_1_187;
   wire n_0_1_188;
   wire n_0_1_189;
   wire n_0_1_190;
   wire n_0_1_191;
   wire n_0_1_192;
   wire n_0_1_193;
   wire n_0_1_194;
   wire n_0_1_195;
   wire n_0_1_196;
   wire n_0_1_197;
   wire n_0_1_198;
   wire n_0_1_199;
   wire n_0_1_200;
   wire n_0_1_201;
   wire n_0_1_202;
   wire n_0_1_203;
   wire n_0_1_204;
   wire n_0_1_205;
   wire n_0_1_206;
   wire n_0_1_207;
   wire n_0_1_208;
   wire n_0_1_209;
   wire n_0_1_210;
   wire n_0_1_211;
   wire n_0_1_212;
   wire n_0_1_213;
   wire n_0_1_214;
   wire n_0_1_215;
   wire n_0_1_216;
   wire n_0_1_217;
   wire n_0_1_218;
   wire n_0_1_219;
   wire n_0_1_220;
   wire n_0_1_221;
   wire n_0_1_222;
   wire n_0_1_223;
   wire [23:0]shiftedToAdd;
   wire n_0_1_224;
   wire n_0_1_225;
   wire n_0_1_226;
   wire n_0_1_227;
   wire n_0_1_228;
   wire n_0_1_229;
   wire n_0_1_230;
   wire n_0_1_231;
   wire n_0_1_232;
   wire n_0_1_233;
   wire n_0_1_234;
   wire n_0_1_235;
   wire n_0_1_236;
   wire n_0_1_237;
   wire n_0_1_238;
   wire n_0_1_239;
   wire n_0_1_240;
   wire n_0_1_241;
   wire n_0_1_242;
   wire n_0_1_243;
   wire n_0_1_244;
   wire n_0_1_245;
   wire n_0_1_246;
   wire n_0_1_247;
   wire n_0_1_248;
   wire n_0_1_249;
   wire n_0_1_250;
   wire n_0_1_251;
   wire n_0_1_252;
   wire n_0_1_253;
   wire n_0_1_254;
   wire n_0_1_255;
   wire n_0_1_256;
   wire n_0_1_257;
   wire n_0_1_258;
   wire n_0_1_259;
   wire n_0_1_260;
   wire n_0_1_261;
   wire n_0_1_262;
   wire n_0_1_263;
   wire n_0_1_264;
   wire n_0_1_265;
   wire n_0_1_266;
   wire n_0_1_267;
   wire n_0_1_268;
   wire n_0_1_269;
   wire n_0_1_270;
   wire n_0_1_271;
   wire n_0_1_272;
   wire n_0_1_273;
   wire n_0_1_274;
   wire n_0_1_275;
   wire n_0_1_276;
   wire n_0_1_277;
   wire n_0_1_278;
   wire n_0_1_279;
   wire n_0_1_280;
   wire n_0_1_281;
   wire n_0_1_282;
   wire n_0_1_283;
   wire n_0_1_284;
   wire n_0_1_285;
   wire n_0_1_286;
   wire n_0_1_287;
   wire n_0_1_288;
   wire n_0_1_289;
   wire n_0_1_290;
   wire n_0_1_291;
   wire n_0_1_292;
   wire n_0_1_293;
   wire n_0_1_294;
   wire n_0_1_295;
   wire n_0_1_296;
   wire n_0_1_297;
   wire n_0_1_298;
   wire n_0_1_299;
   wire n_0_1_300;
   wire n_0_1_301;
   wire n_0_1_302;
   wire n_0_1_303;
   wire n_0_1_304;
   wire n_0_1_305;
   wire n_0_1_306;
   wire n_0_1_307;
   wire n_0_1_308;
   wire n_0_1_309;
   wire n_0_1_310;
   wire n_0_1_311;
   wire n_0_1_312;
   wire n_0_1_313;
   wire n_0_1_314;
   wire n_0_1_315;
   wire n_0_1_316;
   wire n_0_1_317;
   wire n_0_1_318;
   wire n_0_1_319;
   wire n_0_1_320;
   wire n_0_1_321;
   wire n_0_1_322;
   wire n_0_1_323;
   wire n_0_1_324;
   wire n_0_1_325;
   wire n_0_1_326;
   wire n_0_1_327;
   wire n_0_1_328;
   wire n_0_1_329;
   wire n_0_1_330;
   wire n_0_1_331;
   wire n_0_1_332;

   subtractor sub1 (.EA({a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23]}), 
      .EB({b[30], b[29], b[28], b[27], b[26], b[25], b[24], b[23]}), .S2(subsum), 
      .B2(borrow));
   Multiplixer__parameterized0__0_193 Mux2 (.A({a[31], uc_0, a[22], a[21], a[20], 
      a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], a[11], a[10], a[9], 
      a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}), .B({b[31], uc_1, 
      b[22], b[21], b[20], b[19], b[18], b[17], b[16], b[15], b[14], b[13], 
      b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], 
      b[0]}), .Sel(borrow), .Out({outToAdd[24], uc_2, outToAdd[22], outToAdd[21], 
      outToAdd[20], outToAdd[19], outToAdd[18], outToAdd[17], outToAdd[16], 
      outToAdd[15], outToAdd[14], outToAdd[13], outToAdd[12], outToAdd[11], 
      outToAdd[10], outToAdd[9], outToAdd[8], outToAdd[7], outToAdd[6], 
      outToAdd[5], outToAdd[4], outToAdd[3], outToAdd[2], outToAdd[1], 
      outToAdd[0]}));
   Multiplixer__parameterized0 Mux1 (.A({b[31], uc_3, b[22], b[21], b[20], b[19], 
      b[18], b[17], b[16], b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], 
      b[7], b[6], b[5], b[4], b[3], b[2], b[1], b[0]}), .B({a[31], uc_4, a[22], 
      a[21], a[20], a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], 
      a[11], a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}), 
      .Sel(borrow), .Out({outToShift[24], uc_5, outToShift[22], outToShift[21], 
      outToShift[20], outToShift[19], outToShift[18], outToShift[17], 
      outToShift[16], outToShift[15], outToShift[14], outToShift[13], 
      outToShift[12], outToShift[11], outToShift[10], outToShift[9], 
      outToShift[8], outToShift[7], outToShift[6], outToShift[5], outToShift[4], 
      outToShift[3], outToShift[2], outToShift[1], outToShift[0]}));
   CIA_24bit rr (.in1({comA[23], comA[22], comA[21], comA[20], comA[19], 
      comA[18], comA[17], comA[16], comA[15], comA[14], comA[13], comA[12], 
      comA[11], comA[10], comA[9], comA[8], comA[7], comA[6], comA[5], comA[4], 
      comA[3], comA[2], comA[1], shiftedToAdd[0]}), .in2({comB[23], comB[22], 
      comB[21], comB[20], comB[19], comB[18], comB[17], comB[16], comB[15], 
      comB[14], comB[13], comB[12], comB[11], comB[10], comB[9], comB[8], 
      comB[7], comB[6], comB[5], comB[4], comB[3], comB[2], comB[1], outToAdd[0]}), 
      .sum(unNormalizedSum), .carry(carryOfM));
   Multiplixer mux0 (.A({a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23]}), 
      .B({b[30], b[29], b[28], b[27], b[26], b[25], b[24], b[23]}), .Sel(borrow), 
      .Out(ES));
   LZeros lz (.in(unNormalizedSum2), .out(shiftleftamount));
   datapath__0_11 i_0_0 (.p_0({n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_6}), 
      .unNormalizedSum(unNormalizedSum));
   datapath__0_24 i_0_12 (.p_0({n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, 
      n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, uc_7}), 
      .shiftedToAdd(shiftedToAdd));
   datapath__0_27 i_0_15 (.p_0({n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, 
      n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, uc_8}), 
      .outToAdd({uc_9, outToAdd[22], outToAdd[21], outToAdd[20], outToAdd[19], 
      outToAdd[18], outToAdd[17], outToAdd[16], outToAdd[15], outToAdd[14], 
      outToAdd[13], outToAdd[12], outToAdd[11], outToAdd[10], outToAdd[9], 
      outToAdd[8], outToAdd[7], outToAdd[6], outToAdd[5], outToAdd[4], 
      outToAdd[3], outToAdd[2], outToAdd[1], outToAdd[0]}));
   HA_X1 i_0_1_0 (.A(n_0_1_214), .B(ES[0]), .CO(n_0_1_0), .S(n_0_1_14));
   HA_X1 i_0_1_1 (.A(ES[1]), .B(n_0_1_0), .CO(n_0_1_1), .S(n_0_1_15));
   HA_X1 i_0_1_2 (.A(ES[2]), .B(n_0_1_1), .CO(n_0_1_2), .S(n_0_1_16));
   HA_X1 i_0_1_3 (.A(ES[3]), .B(n_0_1_2), .CO(n_0_1_3), .S(n_0_1_17));
   HA_X1 i_0_1_4 (.A(ES[4]), .B(n_0_1_3), .CO(n_0_1_4), .S(n_0_1_18));
   HA_X1 i_0_1_5 (.A(ES[5]), .B(n_0_1_4), .CO(n_0_1_5), .S(n_0_1_19));
   HA_X1 i_0_1_6 (.A(ES[6]), .B(n_0_1_5), .CO(n_0_1_6), .S(n_0_1_20));
   HA_X1 i_0_1_7 (.A(shiftleftamount[0]), .B(ES[0]), .CO(n_0_1_7), .S(n_0_1_21));
   FA_X1 i_0_1_8 (.A(n_0_1_32), .B(ES[1]), .CI(n_0_1_7), .CO(n_0_1_8), .S(
      n_0_1_22));
   FA_X1 i_0_1_9 (.A(n_0_1_31), .B(ES[2]), .CI(n_0_1_8), .CO(n_0_1_9), .S(
      n_0_1_23));
   FA_X1 i_0_1_10 (.A(n_0_1_29), .B(ES[3]), .CI(n_0_1_9), .CO(n_0_1_10), 
      .S(n_0_1_24));
   FA_X1 i_0_1_11 (.A(n_0_1_28), .B(ES[4]), .CI(n_0_1_10), .CO(n_0_1_11), 
      .S(n_0_1_25));
   FA_X1 i_0_1_12 (.A(n_0_1_172), .B(ES[5]), .CI(n_0_1_11), .CO(n_0_1_12), 
      .S(n_0_1_26));
   FA_X1 i_0_1_13 (.A(n_0_1_172), .B(ES[6]), .CI(n_0_1_12), .CO(n_0_1_13), 
      .S(n_0_1_27));
   XNOR2_X1 i_0_1_14 (.A(shiftleftamount[4]), .B(n_0_1_173), .ZN(n_0_1_28));
   NOR2_X1 i_0_1_15 (.A1(n_0_1_173), .A2(n_0_1_30), .ZN(n_0_1_29));
   AOI21_X1 i_0_1_16 (.A(n_0_1_328), .B1(n_0_1_176), .B2(n_0_1_327), .ZN(
      n_0_1_30));
   XNOR2_X1 i_0_1_17 (.A(shiftleftamount[2]), .B(n_0_1_176), .ZN(n_0_1_31));
   XNOR2_X1 i_0_1_18 (.A(n_0_1_326), .B(shiftleftamount[0]), .ZN(n_0_1_32));
   MUX2_X1 i_0_1_19 (.A(n_0_46), .B(outToAdd[1]), .S(n_0_1_223), .Z(comB[1]));
   MUX2_X1 i_0_1_20 (.A(n_0_47), .B(outToAdd[2]), .S(n_0_1_223), .Z(comB[2]));
   MUX2_X1 i_0_1_21 (.A(n_0_48), .B(outToAdd[3]), .S(n_0_1_223), .Z(comB[3]));
   MUX2_X1 i_0_1_22 (.A(n_0_49), .B(outToAdd[4]), .S(n_0_1_223), .Z(comB[4]));
   MUX2_X1 i_0_1_23 (.A(n_0_50), .B(outToAdd[5]), .S(n_0_1_223), .Z(comB[5]));
   MUX2_X1 i_0_1_24 (.A(n_0_51), .B(outToAdd[6]), .S(n_0_1_223), .Z(comB[6]));
   MUX2_X1 i_0_1_25 (.A(n_0_52), .B(outToAdd[7]), .S(n_0_1_223), .Z(comB[7]));
   MUX2_X1 i_0_1_26 (.A(n_0_53), .B(outToAdd[8]), .S(n_0_1_223), .Z(comB[8]));
   MUX2_X1 i_0_1_27 (.A(n_0_54), .B(outToAdd[9]), .S(n_0_1_223), .Z(comB[9]));
   MUX2_X1 i_0_1_28 (.A(n_0_55), .B(outToAdd[10]), .S(n_0_1_223), .Z(comB[10]));
   MUX2_X1 i_0_1_29 (.A(n_0_56), .B(outToAdd[11]), .S(n_0_1_223), .Z(comB[11]));
   MUX2_X1 i_0_1_30 (.A(n_0_57), .B(outToAdd[12]), .S(n_0_1_223), .Z(comB[12]));
   MUX2_X1 i_0_1_31 (.A(n_0_58), .B(outToAdd[13]), .S(n_0_1_223), .Z(comB[13]));
   MUX2_X1 i_0_1_32 (.A(n_0_59), .B(outToAdd[14]), .S(n_0_1_223), .Z(comB[14]));
   MUX2_X1 i_0_1_33 (.A(n_0_60), .B(outToAdd[15]), .S(n_0_1_223), .Z(comB[15]));
   MUX2_X1 i_0_1_34 (.A(n_0_61), .B(outToAdd[16]), .S(n_0_1_223), .Z(comB[16]));
   MUX2_X1 i_0_1_35 (.A(n_0_62), .B(outToAdd[17]), .S(n_0_1_223), .Z(comB[17]));
   MUX2_X1 i_0_1_36 (.A(n_0_63), .B(outToAdd[18]), .S(n_0_1_223), .Z(comB[18]));
   MUX2_X1 i_0_1_37 (.A(n_0_64), .B(outToAdd[19]), .S(n_0_1_223), .Z(comB[19]));
   MUX2_X1 i_0_1_38 (.A(n_0_65), .B(outToAdd[20]), .S(n_0_1_223), .Z(comB[20]));
   MUX2_X1 i_0_1_39 (.A(n_0_66), .B(outToAdd[21]), .S(n_0_1_223), .Z(comB[21]));
   MUX2_X1 i_0_1_40 (.A(n_0_67), .B(outToAdd[22]), .S(n_0_1_223), .Z(comB[22]));
   OR2_X1 i_0_1_41 (.A1(n_0_1_223), .A2(n_0_68), .ZN(comB[23]));
   MUX2_X1 i_0_1_42 (.A(n_0_23), .B(shiftedToAdd[1]), .S(n_0_1_221), .Z(comA[1]));
   MUX2_X1 i_0_1_43 (.A(n_0_24), .B(shiftedToAdd[2]), .S(n_0_1_221), .Z(comA[2]));
   MUX2_X1 i_0_1_44 (.A(n_0_25), .B(shiftedToAdd[3]), .S(n_0_1_221), .Z(comA[3]));
   MUX2_X1 i_0_1_45 (.A(n_0_26), .B(shiftedToAdd[4]), .S(n_0_1_221), .Z(comA[4]));
   MUX2_X1 i_0_1_46 (.A(n_0_27), .B(shiftedToAdd[5]), .S(n_0_1_221), .Z(comA[5]));
   MUX2_X1 i_0_1_47 (.A(n_0_28), .B(shiftedToAdd[6]), .S(n_0_1_221), .Z(comA[6]));
   MUX2_X1 i_0_1_48 (.A(n_0_29), .B(shiftedToAdd[7]), .S(n_0_1_221), .Z(comA[7]));
   MUX2_X1 i_0_1_49 (.A(n_0_30), .B(shiftedToAdd[8]), .S(n_0_1_221), .Z(comA[8]));
   MUX2_X1 i_0_1_50 (.A(n_0_31), .B(shiftedToAdd[9]), .S(n_0_1_221), .Z(comA[9]));
   MUX2_X1 i_0_1_51 (.A(n_0_32), .B(shiftedToAdd[10]), .S(n_0_1_221), .Z(
      comA[10]));
   MUX2_X1 i_0_1_52 (.A(n_0_33), .B(shiftedToAdd[11]), .S(n_0_1_221), .Z(
      comA[11]));
   MUX2_X1 i_0_1_53 (.A(n_0_34), .B(shiftedToAdd[12]), .S(n_0_1_221), .Z(
      comA[12]));
   MUX2_X1 i_0_1_54 (.A(n_0_35), .B(shiftedToAdd[13]), .S(n_0_1_221), .Z(
      comA[13]));
   MUX2_X1 i_0_1_55 (.A(n_0_36), .B(shiftedToAdd[14]), .S(n_0_1_221), .Z(
      comA[14]));
   MUX2_X1 i_0_1_56 (.A(n_0_37), .B(shiftedToAdd[15]), .S(n_0_1_221), .Z(
      comA[15]));
   MUX2_X1 i_0_1_57 (.A(n_0_38), .B(shiftedToAdd[16]), .S(n_0_1_221), .Z(
      comA[16]));
   MUX2_X1 i_0_1_58 (.A(n_0_39), .B(shiftedToAdd[17]), .S(n_0_1_221), .Z(
      comA[17]));
   MUX2_X1 i_0_1_59 (.A(n_0_40), .B(shiftedToAdd[18]), .S(n_0_1_221), .Z(
      comA[18]));
   MUX2_X1 i_0_1_60 (.A(n_0_41), .B(shiftedToAdd[19]), .S(n_0_1_221), .Z(
      comA[19]));
   MUX2_X1 i_0_1_61 (.A(n_0_42), .B(shiftedToAdd[20]), .S(n_0_1_221), .Z(
      comA[20]));
   MUX2_X1 i_0_1_62 (.A(n_0_43), .B(shiftedToAdd[21]), .S(n_0_1_221), .Z(
      comA[21]));
   MUX2_X1 i_0_1_63 (.A(n_0_44), .B(shiftedToAdd[22]), .S(n_0_1_221), .Z(
      comA[22]));
   MUX2_X1 i_0_1_64 (.A(n_0_45), .B(shiftedToAdd[23]), .S(n_0_1_221), .Z(
      comA[23]));
   AND2_X1 i_0_1_65 (.A1(unNormalizedSum2[0]), .A2(n_0_1_33), .ZN(sum[0]));
   NAND2_X1 i_0_1_66 (.A1(n_0_1_220), .A2(n_0_1_172), .ZN(n_0_1_33));
   OAI21_X1 i_0_1_67 (.A(n_0_1_34), .B1(n_0_1_35), .B2(n_0_1_180), .ZN(sum[1]));
   AOI22_X1 i_0_1_68 (.A1(unNormalizedSum[2]), .A2(n_0_1_214), .B1(n_0_1_37), 
      .B2(unNormalizedSum[0]), .ZN(n_0_1_34));
   AOI21_X1 i_0_1_69 (.A(n_0_1_217), .B1(n_0_1_174), .B2(n_0_1_162), .ZN(
      n_0_1_35));
   OAI221_X1 i_0_1_70 (.A(n_0_1_36), .B1(n_0_1_332), .B2(n_0_1_184), .C1(
      n_0_1_39), .C2(n_0_1_161), .ZN(sum[2]));
   AOI22_X1 i_0_1_71 (.A1(n_0_1_181), .A2(n_0_1_37), .B1(unNormalizedSum[3]), 
      .B2(n_0_1_214), .ZN(n_0_1_36));
   NOR3_X1 i_0_1_72 (.A1(n_0_1_177), .A2(n_0_1_175), .A3(n_0_1_137), .ZN(
      n_0_1_37));
   OAI221_X1 i_0_1_73 (.A(n_0_1_38), .B1(n_0_1_39), .B2(n_0_1_137), .C1(
      n_0_1_161), .C2(n_0_1_41), .ZN(sum[3]));
   AOI22_X1 i_0_1_74 (.A1(n_0_1_187), .A2(n_0_1_217), .B1(unNormalizedSum[4]), 
      .B2(n_0_1_214), .ZN(n_0_1_38));
   AOI22_X1 i_0_1_75 (.A1(n_0_1_183), .A2(n_0_1_174), .B1(n_0_1_46), .B2(
      unNormalizedSum[0]), .ZN(n_0_1_39));
   OAI221_X1 i_0_1_76 (.A(n_0_1_40), .B1(n_0_1_41), .B2(n_0_1_137), .C1(
      n_0_1_161), .C2(n_0_1_42), .ZN(sum[4]));
   AOI22_X1 i_0_1_77 (.A1(n_0_1_189), .A2(n_0_1_217), .B1(unNormalizedSum[5]), 
      .B2(n_0_1_214), .ZN(n_0_1_40));
   AOI22_X1 i_0_1_78 (.A1(n_0_1_187), .A2(n_0_1_174), .B1(n_0_1_181), .B2(
      n_0_1_46), .ZN(n_0_1_41));
   AOI221_X1 i_0_1_79 (.A(n_0_1_43), .B1(n_0_1_42), .B2(n_0_1_138), .C1(n_0_1_44), 
      .C2(n_0_1_162), .ZN(sum[5]));
   AOI22_X1 i_0_1_80 (.A1(n_0_1_326), .A2(n_0_1_51), .B1(n_0_1_46), .B2(
      n_0_1_183), .ZN(n_0_1_42));
   OAI22_X1 i_0_1_81 (.A1(n_0_1_332), .A2(n_0_1_191), .B1(n_0_1_215), .B2(
      unNormalizedSum[6]), .ZN(n_0_1_43));
   AOI221_X1 i_0_1_82 (.A(n_0_1_47), .B1(n_0_1_49), .B2(n_0_1_162), .C1(n_0_1_44), 
      .C2(n_0_1_138), .ZN(sum[6]));
   AOI21_X1 i_0_1_83 (.A(n_0_1_45), .B1(n_0_1_46), .B2(n_0_1_187), .ZN(n_0_1_44));
   NOR2_X1 i_0_1_84 (.A1(n_0_1_56), .A2(shiftleftamount[1]), .ZN(n_0_1_45));
   NOR3_X1 i_0_1_85 (.A1(n_0_1_175), .A2(shiftleftamount[2]), .A3(n_0_1_326), 
      .ZN(n_0_1_46));
   OAI22_X1 i_0_1_86 (.A1(n_0_1_332), .A2(n_0_1_192), .B1(n_0_1_215), .B2(
      unNormalizedSum[7]), .ZN(n_0_1_47));
   AOI221_X1 i_0_1_87 (.A(n_0_1_48), .B1(n_0_1_49), .B2(n_0_1_138), .C1(
      n_0_1_162), .C2(n_0_1_54), .ZN(sum[7]));
   OAI22_X1 i_0_1_88 (.A1(n_0_1_332), .A2(n_0_1_197), .B1(n_0_1_215), .B2(
      unNormalizedSum[8]), .ZN(n_0_1_48));
   OAI21_X1 i_0_1_89 (.A(n_0_1_50), .B1(n_0_1_59), .B2(shiftleftamount[1]), 
      .ZN(n_0_1_49));
   NAND2_X1 i_0_1_90 (.A1(n_0_1_52), .A2(shiftleftamount[1]), .ZN(n_0_1_50));
   INV_X1 i_0_1_91 (.A(n_0_1_52), .ZN(n_0_1_51));
   AOI22_X1 i_0_1_92 (.A1(n_0_1_189), .A2(n_0_1_154), .B1(n_0_1_65), .B2(
      unNormalizedSum[0]), .ZN(n_0_1_52));
   AOI221_X1 i_0_1_93 (.A(n_0_1_53), .B1(n_0_1_54), .B2(n_0_1_138), .C1(
      n_0_1_162), .C2(n_0_1_58), .ZN(sum[8]));
   OAI22_X1 i_0_1_94 (.A1(n_0_1_332), .A2(n_0_1_199), .B1(n_0_1_215), .B2(
      unNormalizedSum[9]), .ZN(n_0_1_53));
   OAI21_X1 i_0_1_95 (.A(n_0_1_55), .B1(n_0_1_63), .B2(shiftleftamount[1]), 
      .ZN(n_0_1_54));
   NAND2_X1 i_0_1_96 (.A1(n_0_1_56), .A2(shiftleftamount[1]), .ZN(n_0_1_55));
   AOI22_X1 i_0_1_97 (.A1(n_0_1_191), .A2(n_0_1_154), .B1(n_0_1_181), .B2(
      n_0_1_65), .ZN(n_0_1_56));
   AOI221_X1 i_0_1_98 (.A(n_0_1_57), .B1(n_0_1_58), .B2(n_0_1_138), .C1(
      n_0_1_162), .C2(n_0_1_62), .ZN(sum[9]));
   OAI22_X1 i_0_1_99 (.A1(n_0_1_332), .A2(n_0_1_200), .B1(n_0_1_215), .B2(
      unNormalizedSum[10]), .ZN(n_0_1_57));
   AOI22_X1 i_0_1_100 (.A1(n_0_1_67), .A2(n_0_1_81), .B1(shiftleftamount[1]), 
      .B2(n_0_1_59), .ZN(n_0_1_58));
   INV_X1 i_0_1_101 (.A(n_0_1_60), .ZN(n_0_1_59));
   AOI22_X1 i_0_1_102 (.A1(n_0_1_192), .A2(n_0_1_154), .B1(n_0_1_183), .B2(
      n_0_1_65), .ZN(n_0_1_60));
   AOI221_X1 i_0_1_103 (.A(n_0_1_61), .B1(n_0_1_62), .B2(n_0_1_138), .C1(
      n_0_1_162), .C2(n_0_1_66), .ZN(sum[10]));
   OAI22_X1 i_0_1_104 (.A1(n_0_1_332), .A2(n_0_1_201), .B1(n_0_1_215), .B2(
      unNormalizedSum[11]), .ZN(n_0_1_61));
   AOI22_X1 i_0_1_105 (.A1(n_0_1_70), .A2(n_0_1_81), .B1(shiftleftamount[1]), 
      .B2(n_0_1_63), .ZN(n_0_1_62));
   INV_X1 i_0_1_106 (.A(n_0_1_64), .ZN(n_0_1_63));
   AOI22_X1 i_0_1_107 (.A1(n_0_1_197), .A2(n_0_1_154), .B1(n_0_1_187), .B2(
      n_0_1_65), .ZN(n_0_1_64));
   NOR2_X1 i_0_1_108 (.A1(n_0_1_327), .A2(n_0_1_175), .ZN(n_0_1_65));
   AOI221_X1 i_0_1_109 (.A(n_0_1_68), .B1(n_0_1_66), .B2(n_0_1_138), .C1(
      n_0_1_69), .C2(n_0_1_162), .ZN(sum[11]));
   AOI22_X1 i_0_1_110 (.A1(n_0_1_67), .A2(n_0_1_98), .B1(n_0_1_75), .B2(n_0_1_81), 
      .ZN(n_0_1_66));
   OAI22_X1 i_0_1_111 (.A1(n_0_1_84), .A2(shiftleftamount[2]), .B1(n_0_1_101), 
      .B2(n_0_1_188), .ZN(n_0_1_67));
   OAI22_X1 i_0_1_112 (.A1(n_0_1_332), .A2(n_0_1_202), .B1(n_0_1_215), .B2(
      unNormalizedSum[12]), .ZN(n_0_1_68));
   AOI221_X1 i_0_1_113 (.A(n_0_1_72), .B1(n_0_1_69), .B2(n_0_1_138), .C1(
      n_0_1_73), .C2(n_0_1_162), .ZN(sum[12]));
   AOI22_X1 i_0_1_114 (.A1(n_0_1_81), .A2(n_0_1_78), .B1(n_0_1_70), .B2(n_0_1_98), 
      .ZN(n_0_1_69));
   OAI21_X1 i_0_1_115 (.A(n_0_1_71), .B1(n_0_1_89), .B2(shiftleftamount[2]), 
      .ZN(n_0_1_70));
   NAND3_X1 i_0_1_116 (.A1(n_0_1_328), .A2(n_0_1_191), .A3(shiftleftamount[2]), 
      .ZN(n_0_1_71));
   OAI22_X1 i_0_1_117 (.A1(n_0_1_332), .A2(n_0_1_203), .B1(n_0_1_215), .B2(
      unNormalizedSum[13]), .ZN(n_0_1_72));
   AOI221_X1 i_0_1_118 (.A(n_0_1_76), .B1(n_0_1_162), .B2(n_0_1_77), .C1(
      n_0_1_73), .C2(n_0_1_138), .ZN(sum[13]));
   OAI211_X1 i_0_1_119 (.A(n_0_1_329), .B(n_0_1_74), .C1(n_0_1_75), .C2(
      n_0_1_326), .ZN(n_0_1_73));
   OR2_X1 i_0_1_120 (.A1(n_0_1_82), .A2(shiftleftamount[1]), .ZN(n_0_1_74));
   OAI22_X1 i_0_1_121 (.A1(n_0_1_99), .A2(shiftleftamount[2]), .B1(n_0_1_101), 
      .B2(n_0_1_193), .ZN(n_0_1_75));
   OAI22_X1 i_0_1_122 (.A1(n_0_1_332), .A2(n_0_1_204), .B1(n_0_1_215), .B2(
      unNormalizedSum[14]), .ZN(n_0_1_76));
   AOI221_X1 i_0_1_123 (.A(n_0_1_79), .B1(n_0_1_80), .B2(n_0_1_162), .C1(
      n_0_1_138), .C2(n_0_1_77), .ZN(sum[14]));
   AOI22_X1 i_0_1_124 (.A1(n_0_1_88), .A2(n_0_1_81), .B1(n_0_1_78), .B2(n_0_1_98), 
      .ZN(n_0_1_77));
   OAI22_X1 i_0_1_125 (.A1(shiftleftamount[2]), .A2(n_0_1_105), .B1(n_0_1_101), 
      .B2(n_0_1_196), .ZN(n_0_1_78));
   OAI22_X1 i_0_1_126 (.A1(n_0_1_332), .A2(n_0_1_205), .B1(n_0_1_215), .B2(
      unNormalizedSum[15]), .ZN(n_0_1_79));
   AOI221_X1 i_0_1_127 (.A(n_0_1_86), .B1(n_0_1_80), .B2(n_0_1_138), .C1(
      n_0_1_87), .C2(n_0_1_162), .ZN(sum[15]));
   AOI22_X1 i_0_1_128 (.A1(n_0_1_98), .A2(n_0_1_82), .B1(n_0_1_97), .B2(
      n_0_1_326), .ZN(n_0_1_80));
   NOR2_X1 i_0_1_129 (.A1(shiftleftamount[4]), .A2(shiftleftamount[1]), .ZN(
      n_0_1_81));
   OAI21_X1 i_0_1_130 (.A(n_0_1_83), .B1(n_0_1_84), .B2(n_0_1_327), .ZN(n_0_1_82));
   NAND2_X1 i_0_1_131 (.A1(n_0_1_327), .A2(n_0_1_110), .ZN(n_0_1_83));
   OAI21_X1 i_0_1_132 (.A(n_0_1_85), .B1(unNormalizedSum[0]), .B2(n_0_1_328), 
      .ZN(n_0_1_84));
   OR2_X1 i_0_1_133 (.A1(n_0_1_199), .A2(shiftleftamount[3]), .ZN(n_0_1_85));
   NOR2_X1 i_0_1_134 (.A1(unNormalizedSum2[15]), .A2(n_0_1_220), .ZN(n_0_1_86));
   OAI221_X1 i_0_1_135 (.A(n_0_1_93), .B1(n_0_1_87), .B2(n_0_1_137), .C1(
      n_0_1_95), .C2(n_0_1_161), .ZN(sum[16]));
   AOI22_X1 i_0_1_136 (.A1(n_0_1_326), .A2(n_0_1_104), .B1(n_0_1_98), .B2(
      n_0_1_88), .ZN(n_0_1_87));
   OAI21_X1 i_0_1_137 (.A(n_0_1_92), .B1(n_0_1_89), .B2(n_0_1_327), .ZN(n_0_1_88));
   INV_X1 i_0_1_138 (.A(n_0_1_90), .ZN(n_0_1_89));
   AOI21_X1 i_0_1_139 (.A(n_0_1_91), .B1(n_0_1_180), .B2(shiftleftamount[3]), 
      .ZN(n_0_1_90));
   NOR2_X1 i_0_1_140 (.A1(n_0_1_200), .A2(shiftleftamount[3]), .ZN(n_0_1_91));
   NAND2_X1 i_0_1_141 (.A1(n_0_1_327), .A2(n_0_1_119), .ZN(n_0_1_92));
   AOI22_X1 i_0_1_142 (.A1(unNormalizedSum[16]), .A2(n_0_1_217), .B1(n_0_1_214), 
      .B2(unNormalizedSum[17]), .ZN(n_0_1_93));
   AOI221_X1 i_0_1_143 (.A(n_0_1_94), .B1(n_0_1_102), .B2(n_0_1_162), .C1(
      n_0_1_138), .C2(n_0_1_95), .ZN(sum[17]));
   NOR2_X1 i_0_1_144 (.A1(unNormalizedSum2[17]), .A2(n_0_1_220), .ZN(n_0_1_94));
   OAI21_X1 i_0_1_145 (.A(n_0_1_96), .B1(n_0_1_97), .B2(n_0_1_326), .ZN(n_0_1_95));
   NAND2_X1 i_0_1_146 (.A1(n_0_1_326), .A2(n_0_1_109), .ZN(n_0_1_96));
   OAI22_X1 i_0_1_147 (.A1(n_0_1_127), .A2(n_0_1_123), .B1(n_0_1_99), .B2(
      n_0_1_125), .ZN(n_0_1_97));
   NOR2_X1 i_0_1_148 (.A1(n_0_1_326), .A2(shiftleftamount[4]), .ZN(n_0_1_98));
   OAI21_X1 i_0_1_149 (.A(n_0_1_100), .B1(n_0_1_201), .B2(shiftleftamount[3]), 
      .ZN(n_0_1_99));
   NAND2_X1 i_0_1_150 (.A1(shiftleftamount[3]), .A2(n_0_1_184), .ZN(n_0_1_100));
   NAND2_X1 i_0_1_151 (.A1(n_0_1_328), .A2(shiftleftamount[2]), .ZN(n_0_1_101));
   AOI221_X1 i_0_1_152 (.A(n_0_1_107), .B1(n_0_1_102), .B2(n_0_1_138), .C1(
      n_0_1_108), .C2(n_0_1_162), .ZN(sum[18]));
   OAI21_X1 i_0_1_153 (.A(n_0_1_103), .B1(n_0_1_104), .B2(n_0_1_326), .ZN(
      n_0_1_102));
   OR2_X1 i_0_1_154 (.A1(n_0_1_116), .A2(shiftleftamount[1]), .ZN(n_0_1_103));
   OAI22_X1 i_0_1_155 (.A1(shiftleftamount[2]), .A2(n_0_1_144), .B1(n_0_1_125), 
      .B2(n_0_1_105), .ZN(n_0_1_104));
   OAI21_X1 i_0_1_156 (.A(n_0_1_106), .B1(n_0_1_187), .B2(n_0_1_328), .ZN(
      n_0_1_105));
   OR2_X1 i_0_1_157 (.A1(n_0_1_202), .A2(shiftleftamount[3]), .ZN(n_0_1_106));
   NOR2_X1 i_0_1_158 (.A1(unNormalizedSum2[18]), .A2(n_0_1_220), .ZN(n_0_1_107));
   AOI221_X1 i_0_1_159 (.A(n_0_1_112), .B1(n_0_1_108), .B2(n_0_1_138), .C1(
      n_0_1_114), .C2(n_0_1_162), .ZN(sum[19]));
   MUX2_X1 i_0_1_160 (.A(n_0_1_122), .B(n_0_1_109), .S(shiftleftamount[1]), 
      .Z(n_0_1_108));
   AOI22_X1 i_0_1_161 (.A1(n_0_1_327), .A2(n_0_1_156), .B1(n_0_1_126), .B2(
      n_0_1_110), .ZN(n_0_1_109));
   AOI21_X1 i_0_1_162 (.A(n_0_1_111), .B1(n_0_1_188), .B2(shiftleftamount[3]), 
      .ZN(n_0_1_110));
   NOR2_X1 i_0_1_163 (.A1(n_0_1_203), .A2(shiftleftamount[3]), .ZN(n_0_1_111));
   NOR2_X1 i_0_1_164 (.A1(unNormalizedSum2[19]), .A2(n_0_1_220), .ZN(n_0_1_112));
   OAI221_X1 i_0_1_165 (.A(n_0_1_113), .B1(n_0_1_114), .B2(n_0_1_137), .C1(
      n_0_1_121), .C2(n_0_1_161), .ZN(sum[20]));
   AOI22_X1 i_0_1_166 (.A1(unNormalizedSum[20]), .A2(n_0_1_217), .B1(n_0_1_214), 
      .B2(unNormalizedSum[21]), .ZN(n_0_1_113));
   OAI21_X1 i_0_1_167 (.A(n_0_1_115), .B1(n_0_1_116), .B2(n_0_1_326), .ZN(
      n_0_1_114));
   NAND2_X1 i_0_1_168 (.A1(n_0_1_326), .A2(n_0_1_139), .ZN(n_0_1_115));
   OAI21_X1 i_0_1_169 (.A(n_0_1_117), .B1(n_0_1_118), .B2(n_0_1_125), .ZN(
      n_0_1_116));
   NAND2_X1 i_0_1_170 (.A1(n_0_1_327), .A2(n_0_1_132), .ZN(n_0_1_117));
   INV_X1 i_0_1_171 (.A(n_0_1_119), .ZN(n_0_1_118));
   MUX2_X1 i_0_1_172 (.A(n_0_1_204), .B(n_0_1_191), .S(shiftleftamount[3]), 
      .Z(n_0_1_119));
   OAI21_X1 i_0_1_173 (.A(n_0_1_120), .B1(n_0_1_121), .B2(n_0_1_137), .ZN(
      sum[21]));
   AOI222_X1 i_0_1_174 (.A1(unNormalizedSum[21]), .A2(n_0_1_217), .B1(n_0_1_162), 
      .B2(n_0_1_130), .C1(n_0_1_214), .C2(unNormalizedSum[22]), .ZN(n_0_1_120));
   MUX2_X1 i_0_1_175 (.A(n_0_1_122), .B(n_0_1_151), .S(n_0_1_326), .Z(n_0_1_121));
   AOI21_X1 i_0_1_176 (.A(n_0_1_124), .B1(n_0_1_148), .B2(n_0_1_327), .ZN(
      n_0_1_122));
   NAND2_X1 i_0_1_177 (.A1(n_0_1_329), .A2(n_0_1_327), .ZN(n_0_1_123));
   NOR2_X1 i_0_1_178 (.A1(n_0_1_127), .A2(n_0_1_125), .ZN(n_0_1_124));
   NAND2_X1 i_0_1_179 (.A1(n_0_1_329), .A2(shiftleftamount[2]), .ZN(n_0_1_125));
   NOR2_X1 i_0_1_180 (.A1(n_0_1_327), .A2(shiftleftamount[4]), .ZN(n_0_1_126));
   OAI21_X1 i_0_1_181 (.A(n_0_1_128), .B1(n_0_1_205), .B2(shiftleftamount[3]), 
      .ZN(n_0_1_127));
   NAND2_X1 i_0_1_182 (.A1(shiftleftamount[3]), .A2(n_0_1_193), .ZN(n_0_1_128));
   NAND2_X1 i_0_1_183 (.A1(n_0_1_129), .A2(n_0_1_145), .ZN(sum[22]));
   AOI222_X1 i_0_1_184 (.A1(unNormalizedSum[22]), .A2(n_0_1_217), .B1(n_0_1_138), 
      .B2(n_0_1_130), .C1(n_0_1_214), .C2(unNormalizedSum[23]), .ZN(n_0_1_129));
   AOI221_X1 i_0_1_185 (.A(n_0_1_131), .B1(n_0_1_135), .B2(n_0_1_136), .C1(
      n_0_1_139), .C2(shiftleftamount[1]), .ZN(n_0_1_130));
   NOR2_X1 i_0_1_186 (.A1(n_0_1_146), .A2(n_0_1_132), .ZN(n_0_1_131));
   NAND2_X1 i_0_1_187 (.A1(n_0_1_134), .A2(n_0_1_133), .ZN(n_0_1_132));
   AOI22_X1 i_0_1_188 (.A1(unNormalizedSum[17]), .A2(n_0_1_168), .B1(n_0_1_167), 
      .B2(n_0_16), .ZN(n_0_1_133));
   AOI22_X1 i_0_1_189 (.A1(n_0_1_200), .A2(n_0_1_165), .B1(n_0_1_181), .B2(
      n_0_1_164), .ZN(n_0_1_134));
   AOI22_X1 i_0_1_190 (.A1(n_0_1_204), .A2(n_0_1_165), .B1(n_0_1_191), .B2(
      n_0_1_164), .ZN(n_0_1_135));
   AOI221_X1 i_0_1_191 (.A(n_0_1_177), .B1(n_0_1_168), .B2(unNormalizedSum[21]), 
      .C1(n_0_1_167), .C2(n_0_20), .ZN(n_0_1_136));
   NAND2_X1 i_0_1_192 (.A1(n_0_1_220), .A2(shiftleftamount[0]), .ZN(n_0_1_137));
   NOR2_X1 i_0_1_193 (.A1(n_0_1_330), .A2(n_0_1_325), .ZN(n_0_1_138));
   AOI21_X1 i_0_1_194 (.A(n_0_1_140), .B1(n_0_1_142), .B2(n_0_1_154), .ZN(
      n_0_1_139));
   AOI21_X1 i_0_1_195 (.A(n_0_1_141), .B1(n_0_1_144), .B2(shiftleftamount[2]), 
      .ZN(n_0_1_140));
   AOI221_X1 i_0_1_196 (.A(shiftleftamount[2]), .B1(n_0_1_202), .B2(n_0_1_165), 
      .C1(n_0_1_164), .C2(n_0_1_187), .ZN(n_0_1_141));
   OAI21_X1 i_0_1_197 (.A(n_0_1_143), .B1(n_0_1_331), .B2(n_0_1_317), .ZN(
      n_0_1_142));
   NAND2_X1 i_0_1_198 (.A1(n_0_1_331), .A2(unNormalizedSum[19]), .ZN(n_0_1_143));
   AOI222_X1 i_0_1_199 (.A1(n_0_1_197), .A2(n_0_1_165), .B1(n_0_1_168), .B2(
      unNormalizedSum[15]), .C1(n_0_1_167), .C2(n_0_14), .ZN(n_0_1_144));
   OAI211_X1 i_0_1_200 (.A(n_0_1_147), .B(n_0_1_160), .C1(n_0_1_148), .C2(
      n_0_1_146), .ZN(n_0_1_145));
   NAND2_X1 i_0_1_201 (.A1(n_0_1_326), .A2(shiftleftamount[2]), .ZN(n_0_1_146));
   NAND2_X1 i_0_1_202 (.A1(n_0_1_151), .A2(shiftleftamount[1]), .ZN(n_0_1_147));
   NAND2_X1 i_0_1_203 (.A1(n_0_1_149), .A2(n_0_1_150), .ZN(n_0_1_148));
   AOI22_X1 i_0_1_204 (.A1(n_0_1_201), .A2(n_0_1_165), .B1(n_0_1_183), .B2(
      n_0_1_164), .ZN(n_0_1_149));
   AOI22_X1 i_0_1_205 (.A1(unNormalizedSum[18]), .A2(n_0_1_168), .B1(n_0_1_167), 
      .B2(n_0_17), .ZN(n_0_1_150));
   AOI21_X1 i_0_1_206 (.A(n_0_1_152), .B1(n_0_1_154), .B2(n_0_1_155), .ZN(
      n_0_1_151));
   AOI21_X1 i_0_1_207 (.A(n_0_1_153), .B1(n_0_1_157), .B2(shiftleftamount[2]), 
      .ZN(n_0_1_152));
   AOI221_X1 i_0_1_208 (.A(shiftleftamount[2]), .B1(n_0_1_203), .B2(n_0_1_165), 
      .C1(n_0_1_164), .C2(n_0_1_189), .ZN(n_0_1_153));
   NOR2_X1 i_0_1_209 (.A1(n_0_1_175), .A2(shiftleftamount[2]), .ZN(n_0_1_154));
   MUX2_X1 i_0_1_210 (.A(unNormalizedSum[20]), .B(n_0_19), .S(n_0_1_219), 
      .Z(n_0_1_155));
   INV_X1 i_0_1_211 (.A(n_0_1_157), .ZN(n_0_1_156));
   AOI221_X1 i_0_1_212 (.A(n_0_1_158), .B1(n_0_1_167), .B2(n_0_15), .C1(
      n_0_1_199), .C2(n_0_1_165), .ZN(n_0_1_157));
   INV_X1 i_0_1_213 (.A(n_0_1_159), .ZN(n_0_1_158));
   AOI22_X1 i_0_1_214 (.A1(unNormalizedSum[16]), .A2(n_0_1_168), .B1(n_0_1_164), 
      .B2(unNormalizedSum[0]), .ZN(n_0_1_159));
   AOI21_X1 i_0_1_215 (.A(n_0_1_161), .B1(n_0_1_163), .B2(n_0_1_166), .ZN(
      n_0_1_160));
   NAND2_X1 i_0_1_216 (.A1(n_0_1_325), .A2(n_0_1_220), .ZN(n_0_1_161));
   NOR2_X1 i_0_1_217 (.A1(shiftleftamount[0]), .A2(n_0_1_330), .ZN(n_0_1_162));
   AOI22_X1 i_0_1_218 (.A1(n_0_1_205), .A2(n_0_1_165), .B1(n_0_1_192), .B2(
      n_0_1_164), .ZN(n_0_1_163));
   NOR2_X1 i_0_1_219 (.A1(n_0_1_329), .A2(shiftleftamount[3]), .ZN(n_0_1_164));
   NOR2_X1 i_0_1_220 (.A1(n_0_1_328), .A2(shiftleftamount[4]), .ZN(n_0_1_165));
   AOI221_X1 i_0_1_221 (.A(n_0_1_177), .B1(n_0_1_168), .B2(unNormalizedSum[22]), 
      .C1(n_0_1_167), .C2(n_0_21), .ZN(n_0_1_166));
   NOR2_X1 i_0_1_222 (.A1(n_0_1_331), .A2(n_0_1_175), .ZN(n_0_1_167));
   NOR2_X1 i_0_1_223 (.A1(n_0_1_219), .A2(n_0_1_175), .ZN(n_0_1_168));
   MUX2_X1 i_0_1_224 (.A(n_0_1_14), .B(n_0_1_21), .S(n_0_1_220), .Z(sum[23]));
   MUX2_X1 i_0_1_225 (.A(n_0_1_15), .B(n_0_1_22), .S(n_0_1_220), .Z(sum[24]));
   MUX2_X1 i_0_1_226 (.A(n_0_1_16), .B(n_0_1_23), .S(n_0_1_220), .Z(sum[25]));
   MUX2_X1 i_0_1_227 (.A(n_0_1_17), .B(n_0_1_24), .S(n_0_1_220), .Z(sum[26]));
   MUX2_X1 i_0_1_228 (.A(n_0_1_18), .B(n_0_1_25), .S(n_0_1_220), .Z(sum[27]));
   MUX2_X1 i_0_1_229 (.A(n_0_1_19), .B(n_0_1_26), .S(n_0_1_220), .Z(sum[28]));
   MUX2_X1 i_0_1_230 (.A(n_0_1_20), .B(n_0_1_27), .S(n_0_1_220), .Z(sum[29]));
   XNOR2_X1 i_0_1_231 (.A(ES[7]), .B(n_0_1_169), .ZN(sum[30]));
   OAI21_X1 i_0_1_232 (.A(n_0_1_170), .B1(n_0_1_220), .B2(n_0_1_6), .ZN(
      n_0_1_169));
   NAND2_X1 i_0_1_233 (.A1(n_0_1_220), .A2(n_0_1_171), .ZN(n_0_1_170));
   XNOR2_X1 i_0_1_234 (.A(n_0_1_13), .B(n_0_1_172), .ZN(n_0_1_171));
   NAND2_X1 i_0_1_235 (.A1(n_0_1_174), .A2(n_0_1_325), .ZN(n_0_1_172));
   NOR3_X1 i_0_1_236 (.A1(n_0_1_177), .A2(shiftleftamount[0]), .A3(
      shiftleftamount[3]), .ZN(n_0_1_173));
   NOR2_X1 i_0_1_237 (.A1(n_0_1_177), .A2(n_0_1_175), .ZN(n_0_1_174));
   NAND2_X1 i_0_1_238 (.A1(n_0_1_329), .A2(n_0_1_328), .ZN(n_0_1_175));
   NOR2_X1 i_0_1_239 (.A1(shiftleftamount[1]), .A2(shiftleftamount[0]), .ZN(
      n_0_1_176));
   NAND2_X1 i_0_1_240 (.A1(n_0_1_327), .A2(n_0_1_326), .ZN(n_0_1_177));
   OAI21_X1 i_0_1_241 (.A(n_0_1_179), .B1(n_0_1_178), .B2(carryOfM), .ZN(sum[31]));
   NOR2_X1 i_0_1_242 (.A1(outToShift[24]), .A2(outToAdd[24]), .ZN(n_0_1_178));
   NAND2_X1 i_0_1_243 (.A1(outToShift[24]), .A2(outToAdd[24]), .ZN(n_0_1_179));
   MUX2_X1 i_0_1_244 (.A(unNormalizedSum[1]), .B(unNormalizedSum[0]), .S(
      n_0_1_215), .Z(unNormalizedSum2[0]));
   AOI21_X1 i_0_1_245 (.A(n_0_1_182), .B1(n_0_1_180), .B2(n_0_1_215), .ZN(
      unNormalizedSum2[1]));
   INV_X1 i_0_1_246 (.A(n_0_1_181), .ZN(n_0_1_180));
   MUX2_X1 i_0_1_247 (.A(unNormalizedSum[1]), .B(n_0_0), .S(n_0_1_219), .Z(
      n_0_1_181));
   NOR2_X1 i_0_1_248 (.A1(n_0_1_215), .A2(unNormalizedSum[2]), .ZN(n_0_1_182));
   AOI21_X1 i_0_1_249 (.A(n_0_1_186), .B1(n_0_1_184), .B2(n_0_1_215), .ZN(
      unNormalizedSum2[2]));
   MUX2_X1 i_0_1_250 (.A(unNormalizedSum[2]), .B(n_0_1), .S(n_0_1_219), .Z(
      n_0_1_183));
   AOI21_X1 i_0_1_251 (.A(n_0_1_185), .B1(n_0_1_331), .B2(unNormalizedSum[2]), 
      .ZN(n_0_1_184));
   AND2_X1 i_0_1_252 (.A1(n_0_1), .A2(n_0_1_219), .ZN(n_0_1_185));
   NOR2_X1 i_0_1_253 (.A1(n_0_1_215), .A2(unNormalizedSum[3]), .ZN(n_0_1_186));
   MUX2_X1 i_0_1_254 (.A(unNormalizedSum[4]), .B(n_0_1_187), .S(n_0_1_215), 
      .Z(unNormalizedSum2[3]));
   MUX2_X1 i_0_1_255 (.A(unNormalizedSum[3]), .B(n_0_2), .S(n_0_1_219), .Z(
      n_0_1_187));
   AOI21_X1 i_0_1_256 (.A(n_0_1_190), .B1(n_0_1_188), .B2(n_0_1_215), .ZN(
      unNormalizedSum2[4]));
   INV_X1 i_0_1_257 (.A(n_0_1_189), .ZN(n_0_1_188));
   MUX2_X1 i_0_1_258 (.A(unNormalizedSum[4]), .B(n_0_3), .S(n_0_1_219), .Z(
      n_0_1_189));
   NOR2_X1 i_0_1_259 (.A1(n_0_1_215), .A2(unNormalizedSum[5]), .ZN(n_0_1_190));
   MUX2_X1 i_0_1_260 (.A(unNormalizedSum[6]), .B(n_0_1_191), .S(n_0_1_215), 
      .Z(unNormalizedSum2[5]));
   MUX2_X1 i_0_1_261 (.A(unNormalizedSum[5]), .B(n_0_4), .S(n_0_1_219), .Z(
      n_0_1_191));
   AOI21_X1 i_0_1_262 (.A(n_0_1_195), .B1(n_0_1_193), .B2(n_0_1_215), .ZN(
      unNormalizedSum2[6]));
   MUX2_X1 i_0_1_263 (.A(unNormalizedSum[6]), .B(n_0_5), .S(n_0_1_219), .Z(
      n_0_1_192));
   AOI21_X1 i_0_1_264 (.A(n_0_1_194), .B1(n_0_1_331), .B2(unNormalizedSum[6]), 
      .ZN(n_0_1_193));
   AND2_X1 i_0_1_265 (.A1(n_0_5), .A2(n_0_1_219), .ZN(n_0_1_194));
   NOR2_X1 i_0_1_266 (.A1(n_0_1_215), .A2(unNormalizedSum[7]), .ZN(n_0_1_195));
   AOI21_X1 i_0_1_267 (.A(n_0_1_198), .B1(n_0_1_196), .B2(n_0_1_215), .ZN(
      unNormalizedSum2[7]));
   INV_X1 i_0_1_268 (.A(n_0_1_197), .ZN(n_0_1_196));
   MUX2_X1 i_0_1_269 (.A(unNormalizedSum[7]), .B(n_0_6), .S(n_0_1_219), .Z(
      n_0_1_197));
   NOR2_X1 i_0_1_270 (.A1(n_0_1_215), .A2(unNormalizedSum[8]), .ZN(n_0_1_198));
   MUX2_X1 i_0_1_271 (.A(unNormalizedSum[9]), .B(n_0_1_199), .S(n_0_1_215), 
      .Z(unNormalizedSum2[8]));
   MUX2_X1 i_0_1_272 (.A(unNormalizedSum[8]), .B(n_0_7), .S(n_0_1_219), .Z(
      n_0_1_199));
   MUX2_X1 i_0_1_273 (.A(unNormalizedSum[10]), .B(n_0_1_200), .S(n_0_1_215), 
      .Z(unNormalizedSum2[9]));
   MUX2_X1 i_0_1_274 (.A(unNormalizedSum[9]), .B(n_0_8), .S(n_0_1_219), .Z(
      n_0_1_200));
   MUX2_X1 i_0_1_275 (.A(unNormalizedSum[11]), .B(n_0_1_201), .S(n_0_1_215), 
      .Z(unNormalizedSum2[10]));
   MUX2_X1 i_0_1_276 (.A(unNormalizedSum[10]), .B(n_0_9), .S(n_0_1_219), 
      .Z(n_0_1_201));
   MUX2_X1 i_0_1_277 (.A(unNormalizedSum[12]), .B(n_0_1_202), .S(n_0_1_215), 
      .Z(unNormalizedSum2[11]));
   MUX2_X1 i_0_1_278 (.A(unNormalizedSum[11]), .B(n_0_10), .S(n_0_1_219), 
      .Z(n_0_1_202));
   MUX2_X1 i_0_1_279 (.A(unNormalizedSum[13]), .B(n_0_1_203), .S(n_0_1_215), 
      .Z(unNormalizedSum2[12]));
   MUX2_X1 i_0_1_280 (.A(unNormalizedSum[12]), .B(n_0_11), .S(n_0_1_219), 
      .Z(n_0_1_203));
   MUX2_X1 i_0_1_281 (.A(unNormalizedSum[14]), .B(n_0_1_204), .S(n_0_1_215), 
      .Z(unNormalizedSum2[13]));
   MUX2_X1 i_0_1_282 (.A(unNormalizedSum[13]), .B(n_0_12), .S(n_0_1_219), 
      .Z(n_0_1_204));
   MUX2_X1 i_0_1_283 (.A(unNormalizedSum[15]), .B(n_0_1_205), .S(n_0_1_215), 
      .Z(unNormalizedSum2[14]));
   MUX2_X1 i_0_1_284 (.A(unNormalizedSum[14]), .B(n_0_13), .S(n_0_1_219), 
      .Z(n_0_1_205));
   AOI21_X1 i_0_1_285 (.A(n_0_1_206), .B1(n_0_1_219), .B2(n_0_1_315), .ZN(
      unNormalizedSum2[15]));
   OAI22_X1 i_0_1_286 (.A1(unNormalizedSum[15]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[16]), .ZN(n_0_1_206));
   INV_X1 i_0_1_287 (.A(n_0_1_207), .ZN(unNormalizedSum2[16]));
   OAI222_X1 i_0_1_288 (.A1(unNormalizedSum[16]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[17]), .C1(n_0_1_331), .C2(n_0_15), .ZN(n_0_1_207));
   INV_X1 i_0_1_289 (.A(n_0_1_208), .ZN(unNormalizedSum2[17]));
   OAI222_X1 i_0_1_290 (.A1(unNormalizedSum[17]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[18]), .C1(n_0_1_331), .C2(n_0_16), .ZN(n_0_1_208));
   AOI21_X1 i_0_1_291 (.A(n_0_1_209), .B1(n_0_1_219), .B2(n_0_1_316), .ZN(
      unNormalizedSum2[18]));
   OAI22_X1 i_0_1_292 (.A1(unNormalizedSum[18]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[19]), .ZN(n_0_1_209));
   AOI21_X1 i_0_1_293 (.A(n_0_1_210), .B1(n_0_1_219), .B2(n_0_1_317), .ZN(
      unNormalizedSum2[19]));
   OAI22_X1 i_0_1_294 (.A1(unNormalizedSum[19]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[20]), .ZN(n_0_1_210));
   INV_X1 i_0_1_295 (.A(n_0_1_211), .ZN(unNormalizedSum2[20]));
   OAI222_X1 i_0_1_296 (.A1(unNormalizedSum[20]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[21]), .C1(n_0_1_331), .C2(n_0_19), .ZN(n_0_1_211));
   INV_X1 i_0_1_297 (.A(n_0_1_212), .ZN(unNormalizedSum2[21]));
   OAI222_X1 i_0_1_298 (.A1(unNormalizedSum[21]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[22]), .C1(n_0_1_331), .C2(n_0_20), .ZN(n_0_1_212));
   INV_X1 i_0_1_299 (.A(n_0_1_213), .ZN(unNormalizedSum2[22]));
   OAI222_X1 i_0_1_300 (.A1(unNormalizedSum[22]), .A2(n_0_1_216), .B1(n_0_1_215), 
      .B2(unNormalizedSum[23]), .C1(n_0_1_331), .C2(n_0_21), .ZN(n_0_1_213));
   INV_X1 i_0_1_301 (.A(n_0_1_215), .ZN(n_0_1_214));
   NAND2_X1 i_0_1_302 (.A1(carryOfM), .A2(n_0_1_330), .ZN(n_0_1_215));
   OAI21_X1 i_0_1_303 (.A(n_0_1_218), .B1(n_0_1_216), .B2(n_0_1_324), .ZN(
      unNormalizedSum2[23]));
   XNOR2_X1 i_0_1_304 (.A(carryOfM), .B(n_0_1_330), .ZN(n_0_1_216));
   NOR2_X1 i_0_1_305 (.A1(n_0_1_220), .A2(carryOfM), .ZN(n_0_1_217));
   NAND2_X1 i_0_1_306 (.A1(n_0_22), .A2(n_0_1_219), .ZN(n_0_1_218));
   NOR2_X1 i_0_1_307 (.A1(carryOfM), .A2(n_0_1_330), .ZN(n_0_1_219));
   NAND2_X1 i_0_1_308 (.A1(n_0_1_223), .A2(n_0_1_221), .ZN(n_0_1_220));
   INV_X1 i_0_1_309 (.A(n_0_1_222), .ZN(n_0_1_221));
   NOR2_X1 i_0_1_310 (.A1(n_0_1_319), .A2(outToAdd[24]), .ZN(n_0_1_222));
   NAND2_X1 i_0_1_311 (.A1(n_0_1_319), .A2(outToAdd[24]), .ZN(n_0_1_223));
   OAI22_X1 i_0_1_312 (.A1(n_0_1_298), .A2(n_0_1_228), .B1(n_0_1_224), .B2(
      n_0_1_299), .ZN(shiftedToAdd[0]));
   INV_X1 i_0_1_313 (.A(n_0_1_225), .ZN(n_0_1_224));
   AOI22_X1 i_0_1_314 (.A1(n_0_1_233), .A2(subsum[1]), .B1(n_0_1_226), .B2(
      n_0_1_227), .ZN(n_0_1_225));
   AOI221_X1 i_0_1_315 (.A(subsum[1]), .B1(outToShift[8]), .B2(n_0_1_286), 
      .C1(n_0_1_236), .C2(outToShift[16]), .ZN(n_0_1_226));
   AOI22_X1 i_0_1_316 (.A1(outToShift[0]), .A2(n_0_1_313), .B1(n_0_1_244), 
      .B2(subsum[2]), .ZN(n_0_1_227));
   OAI22_X1 i_0_1_317 (.A1(n_0_1_299), .A2(n_0_1_228), .B1(n_0_1_232), .B2(
      n_0_1_298), .ZN(shiftedToAdd[1]));
   MUX2_X1 i_0_1_318 (.A(n_0_1_229), .B(n_0_1_238), .S(subsum[1]), .Z(n_0_1_228));
   AOI221_X1 i_0_1_319 (.A(n_0_1_230), .B1(n_0_1_313), .B2(outToShift[1]), 
      .C1(subsum[2]), .C2(n_0_1_249), .ZN(n_0_1_229));
   INV_X1 i_0_1_320 (.A(n_0_1_231), .ZN(n_0_1_230));
   AOI22_X1 i_0_1_321 (.A1(outToShift[9]), .A2(n_0_1_286), .B1(n_0_1_236), 
      .B2(outToShift[17]), .ZN(n_0_1_231));
   OAI22_X1 i_0_1_322 (.A1(n_0_1_298), .A2(n_0_1_237), .B1(n_0_1_232), .B2(
      n_0_1_299), .ZN(shiftedToAdd[2]));
   MUX2_X1 i_0_1_323 (.A(n_0_1_233), .B(n_0_1_243), .S(subsum[1]), .Z(n_0_1_232));
   AOI221_X1 i_0_1_324 (.A(n_0_1_234), .B1(n_0_1_286), .B2(outToShift[10]), 
      .C1(subsum[2]), .C2(n_0_1_254), .ZN(n_0_1_233));
   INV_X1 i_0_1_325 (.A(n_0_1_235), .ZN(n_0_1_234));
   AOI22_X1 i_0_1_326 (.A1(outToShift[2]), .A2(n_0_1_313), .B1(n_0_1_236), 
      .B2(outToShift[18]), .ZN(n_0_1_235));
   NOR3_X1 i_0_1_327 (.A1(n_0_1_323), .A2(subsum[3]), .A3(subsum[2]), .ZN(
      n_0_1_236));
   OAI22_X1 i_0_1_328 (.A1(n_0_1_298), .A2(n_0_1_242), .B1(n_0_1_237), .B2(
      n_0_1_299), .ZN(shiftedToAdd[3]));
   MUX2_X1 i_0_1_329 (.A(n_0_1_248), .B(n_0_1_238), .S(n_0_1_321), .Z(n_0_1_237));
   AOI221_X1 i_0_1_330 (.A(n_0_1_239), .B1(n_0_1_313), .B2(outToShift[3]), 
      .C1(outToShift[11]), .C2(n_0_1_286), .ZN(n_0_1_238));
   OAI21_X1 i_0_1_331 (.A(n_0_1_241), .B1(n_0_1_240), .B2(subsum[2]), .ZN(
      n_0_1_239));
   NAND2_X1 i_0_1_332 (.A1(outToShift[19]), .A2(n_0_1_261), .ZN(n_0_1_240));
   NAND2_X1 i_0_1_333 (.A1(subsum[2]), .A2(n_0_1_260), .ZN(n_0_1_241));
   OAI22_X1 i_0_1_334 (.A1(n_0_1_298), .A2(n_0_1_247), .B1(n_0_1_242), .B2(
      n_0_1_299), .ZN(shiftedToAdd[4]));
   MUX2_X1 i_0_1_335 (.A(n_0_1_253), .B(n_0_1_243), .S(n_0_1_321), .Z(n_0_1_242));
   AOI222_X1 i_0_1_336 (.A1(n_0_1_244), .A2(n_0_1_322), .B1(outToShift[8]), 
      .B2(n_0_1_290), .C1(outToShift[16]), .C2(n_0_1_259), .ZN(n_0_1_243));
   NAND2_X1 i_0_1_337 (.A1(n_0_1_246), .A2(n_0_1_245), .ZN(n_0_1_244));
   NAND2_X1 i_0_1_338 (.A1(outToShift[20]), .A2(n_0_1_261), .ZN(n_0_1_245));
   AOI22_X1 i_0_1_339 (.A1(outToShift[4]), .A2(n_0_1_314), .B1(n_0_1_288), 
      .B2(outToShift[12]), .ZN(n_0_1_246));
   OAI22_X1 i_0_1_340 (.A1(n_0_1_298), .A2(n_0_1_252), .B1(n_0_1_247), .B2(
      n_0_1_299), .ZN(shiftedToAdd[5]));
   MUX2_X1 i_0_1_341 (.A(n_0_1_258), .B(n_0_1_248), .S(n_0_1_321), .Z(n_0_1_247));
   AOI222_X1 i_0_1_342 (.A1(n_0_1_249), .A2(n_0_1_322), .B1(outToShift[9]), 
      .B2(n_0_1_290), .C1(outToShift[17]), .C2(n_0_1_259), .ZN(n_0_1_248));
   NAND2_X1 i_0_1_343 (.A1(n_0_1_251), .A2(n_0_1_250), .ZN(n_0_1_249));
   NAND2_X1 i_0_1_344 (.A1(outToShift[21]), .A2(n_0_1_261), .ZN(n_0_1_250));
   AOI22_X1 i_0_1_345 (.A1(outToShift[5]), .A2(n_0_1_314), .B1(n_0_1_288), 
      .B2(outToShift[13]), .ZN(n_0_1_251));
   OAI22_X1 i_0_1_346 (.A1(n_0_1_298), .A2(n_0_1_257), .B1(n_0_1_252), .B2(
      n_0_1_299), .ZN(shiftedToAdd[6]));
   MUX2_X1 i_0_1_347 (.A(n_0_1_263), .B(n_0_1_253), .S(n_0_1_321), .Z(n_0_1_252));
   AOI222_X1 i_0_1_348 (.A1(n_0_1_254), .A2(n_0_1_322), .B1(outToShift[10]), 
      .B2(n_0_1_290), .C1(outToShift[18]), .C2(n_0_1_259), .ZN(n_0_1_253));
   NAND2_X1 i_0_1_349 (.A1(n_0_1_256), .A2(n_0_1_255), .ZN(n_0_1_254));
   NAND2_X1 i_0_1_350 (.A1(outToShift[22]), .A2(n_0_1_261), .ZN(n_0_1_255));
   AOI22_X1 i_0_1_351 (.A1(outToShift[6]), .A2(n_0_1_314), .B1(n_0_1_288), 
      .B2(outToShift[14]), .ZN(n_0_1_256));
   OAI22_X1 i_0_1_352 (.A1(n_0_1_298), .A2(n_0_1_262), .B1(n_0_1_257), .B2(
      n_0_1_299), .ZN(shiftedToAdd[7]));
   MUX2_X1 i_0_1_353 (.A(n_0_1_265), .B(n_0_1_258), .S(n_0_1_321), .Z(n_0_1_257));
   AOI222_X1 i_0_1_354 (.A1(n_0_1_322), .A2(n_0_1_260), .B1(n_0_1_259), .B2(
      outToShift[19]), .C1(outToShift[11]), .C2(n_0_1_290), .ZN(n_0_1_258));
   NOR2_X1 i_0_1_355 (.A1(n_0_1_322), .A2(n_0_1_287), .ZN(n_0_1_259));
   AOI22_X1 i_0_1_356 (.A1(n_0_1_318), .A2(n_0_1_314), .B1(n_0_1_283), .B2(
      subsum[3]), .ZN(n_0_1_260));
   NOR2_X1 i_0_1_357 (.A1(n_0_1_323), .A2(subsum[3]), .ZN(n_0_1_261));
   OAI22_X1 i_0_1_358 (.A1(n_0_1_262), .A2(n_0_1_299), .B1(n_0_1_264), .B2(
      n_0_1_298), .ZN(shiftedToAdd[8]));
   MUX2_X1 i_0_1_359 (.A(n_0_1_267), .B(n_0_1_263), .S(n_0_1_321), .Z(n_0_1_262));
   AOI222_X1 i_0_1_360 (.A1(n_0_1_278), .A2(n_0_1_288), .B1(n_0_1_313), .B2(
      outToShift[8]), .C1(n_0_1_290), .C2(outToShift[12]), .ZN(n_0_1_263));
   OAI22_X1 i_0_1_361 (.A1(n_0_1_266), .A2(n_0_1_298), .B1(n_0_1_299), .B2(
      n_0_1_264), .ZN(shiftedToAdd[9]));
   MUX2_X1 i_0_1_362 (.A(n_0_1_269), .B(n_0_1_265), .S(n_0_1_321), .Z(n_0_1_264));
   AOI222_X1 i_0_1_363 (.A1(n_0_1_294), .A2(n_0_1_288), .B1(n_0_1_290), .B2(
      outToShift[13]), .C1(n_0_1_313), .C2(outToShift[9]), .ZN(n_0_1_265));
   OAI22_X1 i_0_1_364 (.A1(n_0_1_266), .A2(n_0_1_299), .B1(n_0_1_268), .B2(
      n_0_1_298), .ZN(shiftedToAdd[10]));
   MUX2_X1 i_0_1_365 (.A(n_0_1_267), .B(n_0_1_273), .S(subsum[1]), .Z(n_0_1_266));
   AOI222_X1 i_0_1_366 (.A1(n_0_1_296), .A2(n_0_1_288), .B1(n_0_1_290), .B2(
      outToShift[14]), .C1(n_0_1_313), .C2(outToShift[10]), .ZN(n_0_1_267));
   OAI22_X1 i_0_1_367 (.A1(n_0_1_298), .A2(n_0_1_272), .B1(n_0_1_268), .B2(
      n_0_1_299), .ZN(shiftedToAdd[11]));
   MUX2_X1 i_0_1_368 (.A(n_0_1_269), .B(n_0_1_276), .S(subsum[1]), .Z(n_0_1_268));
   OAI211_X1 i_0_1_369 (.A(n_0_1_323), .B(n_0_1_270), .C1(n_0_1_271), .C2(
      subsum[3]), .ZN(n_0_1_269));
   NAND2_X1 i_0_1_370 (.A1(subsum[3]), .A2(n_0_1_304), .ZN(n_0_1_270));
   MUX2_X1 i_0_1_371 (.A(outToShift[11]), .B(outToShift[15]), .S(subsum[2]), 
      .Z(n_0_1_271));
   OAI22_X1 i_0_1_372 (.A1(n_0_1_272), .A2(n_0_1_299), .B1(n_0_1_274), .B2(
      n_0_1_298), .ZN(shiftedToAdd[12]));
   MUX2_X1 i_0_1_373 (.A(n_0_1_280), .B(n_0_1_273), .S(n_0_1_321), .Z(n_0_1_272));
   AOI222_X1 i_0_1_374 (.A1(outToShift[12]), .A2(n_0_1_313), .B1(n_0_1_290), 
      .B2(outToShift[16]), .C1(outToShift[20]), .C2(n_0_1_286), .ZN(n_0_1_273));
   OAI22_X1 i_0_1_375 (.A1(n_0_1_277), .A2(n_0_1_298), .B1(n_0_1_299), .B2(
      n_0_1_274), .ZN(shiftedToAdd[13]));
   OAI21_X1 i_0_1_376 (.A(n_0_1_275), .B1(n_0_1_282), .B2(n_0_1_321), .ZN(
      n_0_1_274));
   NAND2_X1 i_0_1_377 (.A1(n_0_1_321), .A2(n_0_1_276), .ZN(n_0_1_275));
   AOI222_X1 i_0_1_378 (.A1(outToShift[13]), .A2(n_0_1_313), .B1(n_0_1_290), 
      .B2(outToShift[17]), .C1(outToShift[21]), .C2(n_0_1_286), .ZN(n_0_1_276));
   OAI22_X1 i_0_1_379 (.A1(n_0_1_277), .A2(n_0_1_299), .B1(n_0_1_281), .B2(
      n_0_1_298), .ZN(shiftedToAdd[14]));
   AOI21_X1 i_0_1_380 (.A(n_0_1_279), .B1(n_0_1_278), .B2(n_0_1_293), .ZN(
      n_0_1_277));
   MUX2_X1 i_0_1_381 (.A(outToShift[16]), .B(outToShift[20]), .S(subsum[2]), 
      .Z(n_0_1_278));
   NOR2_X1 i_0_1_382 (.A1(n_0_1_280), .A2(subsum[1]), .ZN(n_0_1_279));
   AOI222_X1 i_0_1_383 (.A1(outToShift[14]), .A2(n_0_1_313), .B1(n_0_1_290), 
      .B2(outToShift[18]), .C1(outToShift[22]), .C2(n_0_1_286), .ZN(n_0_1_280));
   OAI22_X1 i_0_1_384 (.A1(n_0_1_281), .A2(n_0_1_299), .B1(n_0_1_298), .B2(
      n_0_1_289), .ZN(shiftedToAdd[15]));
   AOI22_X1 i_0_1_385 (.A1(n_0_1_282), .A2(n_0_1_321), .B1(n_0_1_293), .B2(
      n_0_1_294), .ZN(n_0_1_281));
   OAI211_X1 i_0_1_386 (.A(n_0_1_285), .B(n_0_1_284), .C1(n_0_1_283), .C2(
      subsum[2]), .ZN(n_0_1_282));
   NAND2_X1 i_0_1_387 (.A1(n_0_1_323), .A2(outToShift[15]), .ZN(n_0_1_283));
   NAND3_X1 i_0_1_388 (.A1(subsum[2]), .A2(outToShift[19]), .A3(n_0_1_314), 
      .ZN(n_0_1_284));
   INV_X1 i_0_1_389 (.A(n_0_1_286), .ZN(n_0_1_285));
   NOR2_X1 i_0_1_390 (.A1(n_0_1_287), .A2(subsum[2]), .ZN(n_0_1_286));
   INV_X1 i_0_1_391 (.A(n_0_1_288), .ZN(n_0_1_287));
   AND2_X1 i_0_1_392 (.A1(n_0_1_323), .A2(subsum[3]), .ZN(n_0_1_288));
   OAI22_X1 i_0_1_393 (.A1(n_0_1_298), .A2(n_0_1_292), .B1(n_0_1_289), .B2(
      n_0_1_299), .ZN(shiftedToAdd[16]));
   AOI22_X1 i_0_1_394 (.A1(n_0_1_306), .A2(n_0_1_290), .B1(n_0_1_291), .B2(
      n_0_1_313), .ZN(n_0_1_289));
   NOR3_X1 i_0_1_395 (.A1(n_0_1_322), .A2(subsum[3]), .A3(subsum[4]), .ZN(
      n_0_1_290));
   MUX2_X1 i_0_1_396 (.A(outToShift[16]), .B(outToShift[18]), .S(subsum[1]), 
      .Z(n_0_1_291));
   OAI22_X1 i_0_1_397 (.A1(n_0_1_298), .A2(n_0_1_295), .B1(n_0_1_292), .B2(
      n_0_1_299), .ZN(shiftedToAdd[17]));
   AOI22_X1 i_0_1_398 (.A1(n_0_1_302), .A2(n_0_1_294), .B1(n_0_1_293), .B2(
      n_0_1_303), .ZN(n_0_1_292));
   NOR3_X1 i_0_1_399 (.A1(n_0_1_321), .A2(subsum[3]), .A3(subsum[4]), .ZN(
      n_0_1_293));
   MUX2_X1 i_0_1_400 (.A(outToShift[17]), .B(outToShift[21]), .S(subsum[2]), 
      .Z(n_0_1_294));
   OAI22_X1 i_0_1_401 (.A1(n_0_1_300), .A2(n_0_1_298), .B1(n_0_1_295), .B2(
      n_0_1_299), .ZN(shiftedToAdd[18]));
   AOI22_X1 i_0_1_402 (.A1(n_0_1_302), .A2(n_0_1_296), .B1(n_0_1_301), .B2(
      outToShift[20]), .ZN(n_0_1_295));
   MUX2_X1 i_0_1_403 (.A(outToShift[18]), .B(outToShift[22]), .S(subsum[2]), 
      .Z(n_0_1_296));
   OAI22_X1 i_0_1_404 (.A1(n_0_1_300), .A2(n_0_1_299), .B1(n_0_1_298), .B2(
      n_0_1_297), .ZN(shiftedToAdd[19]));
   NAND2_X1 i_0_1_405 (.A1(n_0_1_306), .A2(n_0_1_313), .ZN(n_0_1_297));
   NAND2_X1 i_0_1_406 (.A1(subsum[0]), .A2(n_0_1_312), .ZN(n_0_1_298));
   NAND2_X1 i_0_1_407 (.A1(n_0_1_312), .A2(n_0_1_320), .ZN(n_0_1_299));
   AOI22_X1 i_0_1_408 (.A1(outToShift[21]), .A2(n_0_1_301), .B1(n_0_1_302), 
      .B2(n_0_1_303), .ZN(n_0_1_300));
   AND2_X1 i_0_1_409 (.A1(subsum[1]), .A2(n_0_1_313), .ZN(n_0_1_301));
   NOR3_X1 i_0_1_410 (.A1(subsum[4]), .A2(subsum[3]), .A3(subsum[1]), .ZN(
      n_0_1_302));
   INV_X1 i_0_1_411 (.A(n_0_1_304), .ZN(n_0_1_303));
   NOR2_X1 i_0_1_412 (.A1(subsum[2]), .A2(outToShift[19]), .ZN(n_0_1_304));
   AOI21_X1 i_0_1_413 (.A(n_0_1_311), .B1(n_0_1_307), .B2(n_0_1_305), .ZN(
      shiftedToAdd[20]));
   NAND2_X1 i_0_1_414 (.A1(n_0_1_320), .A2(n_0_1_306), .ZN(n_0_1_305));
   MUX2_X1 i_0_1_415 (.A(outToShift[20]), .B(outToShift[22]), .S(subsum[1]), 
      .Z(n_0_1_306));
   OAI21_X1 i_0_1_416 (.A(subsum[0]), .B1(outToShift[21]), .B2(subsum[1]), 
      .ZN(n_0_1_307));
   AOI21_X1 i_0_1_417 (.A(n_0_1_311), .B1(n_0_1_309), .B2(n_0_1_308), .ZN(
      shiftedToAdd[21]));
   NAND3_X1 i_0_1_418 (.A1(n_0_1_321), .A2(subsum[0]), .A3(outToShift[22]), 
      .ZN(n_0_1_308));
   OAI21_X1 i_0_1_419 (.A(n_0_1_320), .B1(outToShift[21]), .B2(subsum[1]), 
      .ZN(n_0_1_309));
   NOR3_X1 i_0_1_420 (.A1(n_0_1_311), .A2(n_0_1_310), .A3(subsum[1]), .ZN(
      shiftedToAdd[22]));
   NOR2_X1 i_0_1_421 (.A1(subsum[0]), .A2(outToShift[22]), .ZN(n_0_1_310));
   NOR3_X1 i_0_1_422 (.A1(n_0_1_311), .A2(subsum[0]), .A3(subsum[1]), .ZN(
      shiftedToAdd[23]));
   NAND2_X1 i_0_1_423 (.A1(n_0_1_313), .A2(n_0_1_312), .ZN(n_0_1_311));
   NOR3_X1 i_0_1_424 (.A1(subsum[7]), .A2(subsum[6]), .A3(subsum[5]), .ZN(
      n_0_1_312));
   NOR3_X1 i_0_1_425 (.A1(subsum[4]), .A2(subsum[3]), .A3(subsum[2]), .ZN(
      n_0_1_313));
   NOR2_X1 i_0_1_426 (.A1(subsum[4]), .A2(subsum[3]), .ZN(n_0_1_314));
   INV_X1 i_0_1_427 (.A(n_0_14), .ZN(n_0_1_315));
   INV_X1 i_0_1_428 (.A(n_0_17), .ZN(n_0_1_316));
   INV_X1 i_0_1_429 (.A(n_0_18), .ZN(n_0_1_317));
   INV_X1 i_0_1_430 (.A(outToShift[7]), .ZN(n_0_1_318));
   INV_X1 i_0_1_431 (.A(outToShift[24]), .ZN(n_0_1_319));
   INV_X1 i_0_1_432 (.A(subsum[0]), .ZN(n_0_1_320));
   INV_X1 i_0_1_433 (.A(subsum[1]), .ZN(n_0_1_321));
   INV_X1 i_0_1_434 (.A(subsum[2]), .ZN(n_0_1_322));
   INV_X1 i_0_1_435 (.A(subsum[4]), .ZN(n_0_1_323));
   INV_X1 i_0_1_436 (.A(unNormalizedSum[23]), .ZN(n_0_1_324));
   INV_X1 i_0_1_437 (.A(shiftleftamount[0]), .ZN(n_0_1_325));
   INV_X1 i_0_1_438 (.A(shiftleftamount[1]), .ZN(n_0_1_326));
   INV_X1 i_0_1_439 (.A(shiftleftamount[2]), .ZN(n_0_1_327));
   INV_X1 i_0_1_440 (.A(shiftleftamount[3]), .ZN(n_0_1_328));
   INV_X1 i_0_1_441 (.A(shiftleftamount[4]), .ZN(n_0_1_329));
   INV_X1 i_0_1_442 (.A(n_0_1_220), .ZN(n_0_1_330));
   INV_X1 i_0_1_443 (.A(n_0_1_219), .ZN(n_0_1_331));
   INV_X1 i_0_1_444 (.A(n_0_1_217), .ZN(n_0_1_332));
endmodule
